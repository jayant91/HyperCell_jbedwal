module ALU(
    input [31:0] io_inOp1,
    input [31:0] io_inOp2,
    output[31:0] io_out,
    input [4:0] io_opCode,
    input  io_inOp1Valid,
    input  io_inOp2Valid,
    output io_outValid
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire[31:0] T196;
  wire[63:0] T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire[63:0] T139;
  wire[63:0] T140;
  wire[63:0] T141;
  wire[63:0] T142;
  wire[63:0] T143;
  wire[63:0] T144;
  wire[63:0] T145;
  wire[63:0] T146;
  wire[63:0] T147;
  wire[63:0] T148;
  wire[63:0] T149;
  wire[63:0] T150;
  wire[63:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[63:0] T154;
  wire[63:0] T155;
  wire[63:0] T156;
  wire[63:0] T157;
  wire[63:0] T158;
  wire[63:0] T197;
  wire[31:0] T159;
  wire[31:0] T160;
  wire[31:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  wire[63:0] T165;
  wire[63:0] T198;
  wire[31:0] T166;
  wire[63:0] T199;
  wire[31:0] T167;
  wire[63:0] T200;
  wire[31:0] T168;
  wire[63:0] T201;
  wire[31:0] T169;
  wire[63:0] T202;
  wire[31:0] T170;
  wire[63:0] T203;
  wire[31:0] T171;
  wire[63:0] T204;
  wire[31:0] T172;
  wire[31:0] tempInS;
  wire[31:0] T205;
  wire[32:0] T173;
  wire[32:0] T174;
  wire[32:0] T175;
  wire[31:0] T206;
  wire T207;
  wire[63:0] T208;
  wire[31:0] T176;
  wire[31:0] temp2;
  wire[31:0] T209;
  wire[94:0] T177;
  wire[94:0] T178;
  wire[94:0] T179;
  wire[5:0] T180;
  wire[5:0] T181;
  wire[94:0] T210;
  wire[31:0] T182;
  wire[5:0] T183;
  wire[5:0] T184;
  wire[31:0] temp1;
  wire[31:0] T211;
  wire[94:0] T185;
  wire[94:0] T212;
  wire[31:0] T186;
  wire[31:0] T187;
  wire[5:0] T188;
  wire[94:0] T189;
  wire[5:0] T190;
  wire[63:0] T213;
  wire[31:0] T191;
  wire[63:0] T214;
  wire[31:0] T192;
  wire T193;
  wire[63:0] T215;
  wire[31:0] T194;
  wire T195;


  assign io_outValid = T0;
  assign T0 = T133 ? 1'h0 : T1;
  assign T1 = T127 ? 1'h1 : T2;
  assign T2 = T125 ? 1'h0 : T3;
  assign T3 = T119 ? 1'h1 : T4;
  assign T4 = T117 ? 1'h0 : T5;
  assign T5 = T111 ? 1'h1 : T6;
  assign T6 = T109 ? 1'h0 : T7;
  assign T7 = T103 ? 1'h1 : T8;
  assign T8 = T101 ? 1'h0 : T9;
  assign T9 = T95 ? 1'h1 : T10;
  assign T10 = T93 ? 1'h0 : T11;
  assign T11 = T87 ? 1'h1 : T12;
  assign T12 = T85 ? 1'h0 : T13;
  assign T13 = T79 ? 1'h1 : T14;
  assign T14 = T77 ? 1'h0 : T15;
  assign T15 = T72 ? 1'h1 : T16;
  assign T16 = T70 ? 1'h0 : T17;
  assign T17 = T64 ? 1'h1 : T18;
  assign T18 = T62 ? 1'h0 : T19;
  assign T19 = T56 ? 1'h1 : T20;
  assign T20 = T54 ? 1'h0 : T21;
  assign T21 = T48 ? 1'h1 : T22;
  assign T22 = T46 ? 1'h0 : T23;
  assign T23 = T40 ? 1'h1 : T24;
  assign T24 = T38 ? 1'h0 : T25;
  assign T25 = T33 ? 1'h1 : T26;
  assign T26 = T31 ? 1'h0 : T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = T30 & T29;
  assign T29 = io_inOp1Valid & io_inOp2Valid;
  assign T30 = io_opCode == 5'h0;
  assign T31 = T30 & T32;
  assign T32 = T29 ^ 1'h1;
  assign T33 = T35 & T34;
  assign T34 = io_inOp1Valid & io_inOp2Valid;
  assign T35 = T37 & T36;
  assign T36 = io_opCode == 5'h1;
  assign T37 = T30 ^ 1'h1;
  assign T38 = T35 & T39;
  assign T39 = T34 ^ 1'h1;
  assign T40 = T42 & T41;
  assign T41 = io_inOp1Valid & io_inOp2Valid;
  assign T42 = T44 & T43;
  assign T43 = io_opCode == 5'h2;
  assign T44 = T45 ^ 1'h1;
  assign T45 = T30 | T36;
  assign T46 = T42 & T47;
  assign T47 = T41 ^ 1'h1;
  assign T48 = T50 & T49;
  assign T49 = io_inOp1Valid & io_inOp2Valid;
  assign T50 = T52 & T51;
  assign T51 = io_opCode == 5'h3;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T45 | T43;
  assign T54 = T50 & T55;
  assign T55 = T49 ^ 1'h1;
  assign T56 = T58 & T57;
  assign T57 = io_inOp1Valid & io_inOp2Valid;
  assign T58 = T60 & T59;
  assign T59 = io_opCode == 5'h4;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T53 | T51;
  assign T62 = T58 & T63;
  assign T63 = T57 ^ 1'h1;
  assign T64 = T66 & T65;
  assign T65 = io_inOp1Valid & io_inOp2Valid;
  assign T66 = T68 & T67;
  assign T67 = io_opCode == 5'h5;
  assign T68 = T69 ^ 1'h1;
  assign T69 = T61 | T59;
  assign T70 = T66 & T71;
  assign T71 = T65 ^ 1'h1;
  assign T72 = T73 & io_inOp1Valid;
  assign T73 = T75 & T74;
  assign T74 = io_opCode == 5'h6;
  assign T75 = T76 ^ 1'h1;
  assign T76 = T69 | T67;
  assign T77 = T73 & T78;
  assign T78 = io_inOp1Valid ^ 1'h1;
  assign T79 = T81 & T80;
  assign T80 = io_inOp1Valid & io_inOp2Valid;
  assign T81 = T83 & T82;
  assign T82 = io_opCode == 5'h7;
  assign T83 = T84 ^ 1'h1;
  assign T84 = T76 | T74;
  assign T85 = T81 & T86;
  assign T86 = T80 ^ 1'h1;
  assign T87 = T89 & T88;
  assign T88 = io_inOp1Valid & io_inOp2Valid;
  assign T89 = T91 & T90;
  assign T90 = io_opCode == 5'h8;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T84 | T82;
  assign T93 = T89 & T94;
  assign T94 = T88 ^ 1'h1;
  assign T95 = T97 & T96;
  assign T96 = io_inOp1Valid & io_inOp2Valid;
  assign T97 = T99 & T98;
  assign T98 = io_opCode == 5'h9;
  assign T99 = T100 ^ 1'h1;
  assign T100 = T92 | T90;
  assign T101 = T97 & T102;
  assign T102 = T96 ^ 1'h1;
  assign T103 = T105 & T104;
  assign T104 = io_inOp1Valid & io_inOp2Valid;
  assign T105 = T107 & T106;
  assign T106 = io_opCode == 5'ha;
  assign T107 = T108 ^ 1'h1;
  assign T108 = T100 | T98;
  assign T109 = T105 & T110;
  assign T110 = T104 ^ 1'h1;
  assign T111 = T113 & T112;
  assign T112 = io_inOp1Valid & io_inOp2Valid;
  assign T113 = T115 & T114;
  assign T114 = io_opCode == 5'hb;
  assign T115 = T116 ^ 1'h1;
  assign T116 = T108 | T106;
  assign T117 = T113 & T118;
  assign T118 = T112 ^ 1'h1;
  assign T119 = T121 & T120;
  assign T120 = io_inOp1Valid & io_inOp2Valid;
  assign T121 = T123 & T122;
  assign T122 = io_opCode == 5'hc;
  assign T123 = T124 ^ 1'h1;
  assign T124 = T116 | T114;
  assign T125 = T121 & T126;
  assign T126 = T120 ^ 1'h1;
  assign T127 = T129 & T128;
  assign T128 = io_inOp1Valid & io_inOp2Valid;
  assign T129 = T131 & T130;
  assign T130 = io_opCode == 5'hd;
  assign T131 = T132 ^ 1'h1;
  assign T132 = T124 | T122;
  assign T133 = T129 & T134;
  assign T134 = T128 ^ 1'h1;
  assign io_out = T196;
  assign T196 = T135[5'h1f:1'h0];
  assign T135 = T133 ? 64'h0 : T136;
  assign T136 = T127 ? T215 : T137;
  assign T137 = T125 ? 64'h0 : T138;
  assign T138 = T119 ? T214 : T139;
  assign T139 = T117 ? 64'h0 : T140;
  assign T140 = T111 ? T213 : T141;
  assign T141 = T109 ? 64'h0 : T142;
  assign T142 = T103 ? T208 : T143;
  assign T143 = T101 ? 64'h0 : T144;
  assign T144 = T95 ? T204 : T145;
  assign T145 = T93 ? 64'h0 : T146;
  assign T146 = T87 ? T203 : T147;
  assign T147 = T85 ? 64'h0 : T148;
  assign T148 = T79 ? T202 : T149;
  assign T149 = T77 ? 64'h0 : T150;
  assign T150 = T72 ? T201 : T151;
  assign T151 = T70 ? 64'h0 : T152;
  assign T152 = T64 ? T200 : T153;
  assign T153 = T62 ? 64'h0 : T154;
  assign T154 = T56 ? T199 : T155;
  assign T155 = T54 ? 64'h0 : T156;
  assign T156 = T48 ? T198 : T157;
  assign T157 = T46 ? 64'h0 : T158;
  assign T158 = T40 ? T165 : T197;
  assign T197 = {32'h0, T159};
  assign T159 = T38 ? 32'h0 : T160;
  assign T160 = T33 ? T164 : T161;
  assign T161 = T31 ? 32'h0 : T162;
  assign T162 = T28 ? T163 : 32'h0;
  assign T163 = io_inOp1 + io_inOp2;
  assign T164 = io_inOp1 - io_inOp2;
  assign T165 = io_inOp1 * io_inOp2;
  assign T198 = {32'h0, T166};
  assign T166 = io_inOp1 & io_inOp2;
  assign T199 = {32'h0, T167};
  assign T167 = io_inOp1 | io_inOp2;
  assign T200 = {32'h0, T168};
  assign T168 = io_inOp1 ^ io_inOp2;
  assign T201 = {32'h0, T169};
  assign T169 = ~ io_inOp1;
  assign T202 = {32'h0, T170};
  assign T170 = io_inOp1 << io_inOp2;
  assign T203 = {32'h0, T171};
  assign T171 = io_inOp1 >> io_inOp2;
  assign T204 = {T206, T172};
  assign T172 = $signed(tempInS) >>> io_inOp2;
  assign tempInS = T205;
  assign T205 = T173[5'h1f:1'h0];
  assign T173 = T95 ? T174 : 33'h0;
  assign T174 = T175;
  assign T175 = {1'h0, io_inOp1};
  assign T206 = T207 ? 32'hffffffff : 32'h0;
  assign T207 = T172[5'h1f:5'h1f];
  assign T208 = {32'h0, T176};
  assign T176 = temp1 + temp2;
  assign temp2 = T209;
  assign T209 = T177[5'h1f:1'h0];
  assign T177 = T111 ? T210 : T178;
  assign T178 = T103 ? T179 : 95'h0;
  assign T179 = io_inOp1 << T180;
  assign T180 = 6'h20 - T181;
  assign T181 = io_inOp2 % 6'h20;
  assign T210 = {63'h0, T182};
  assign T182 = io_inOp1 >> T183;
  assign T183 = 6'h20 - T184;
  assign T184 = io_inOp2 % 6'h20;
  assign temp1 = T211;
  assign T211 = T185[5'h1f:1'h0];
  assign T185 = T111 ? T189 : T212;
  assign T212 = {63'h0, T186};
  assign T186 = T103 ? T187 : 32'h0;
  assign T187 = io_inOp1 >> T188;
  assign T188 = io_inOp2 % 6'h20;
  assign T189 = io_inOp1 << T190;
  assign T190 = io_inOp2 % 6'h20;
  assign T213 = {32'h0, T191};
  assign T191 = temp1 + temp2;
  assign T214 = {32'h0, T192};
  assign T192 = T193 ? io_inOp1 : io_inOp2;
  assign T193 = io_inOp2 <= io_inOp1;
  assign T215 = {32'h0, T194};
  assign T194 = T195 ? io_inOp1 : io_inOp2;
  assign T195 = io_inOp1 <= io_inOp2;
endmodule

module FifoCU(input clk, input reset,
    input [31:0] io_enqData,
    output[31:0] io_deqData,
    output io_enqRdy,
    input [3:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [3:0] io_deqReg,
    output io_enqRdyOut
);

  wire T0;
  wire T1;
  reg  isFull;
  wire T37;
  wire isFullNext;
  wire T2;
  wire T3;
  wire doDeq;
  wire T4;
  wire T5;
  reg  deqPtr;
  wire T38;
  wire T6;
  wire deqPtrInc;
  wire T7;
  wire enqPtrInc;
  wire T8;
  reg  enqPtr;
  wire T39;
  wire T9;
  wire doEnq;
  wire T10;
  wire T11;
  wire T12;
  wire deqCombined;
  wire[3:0] deqCond;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire isEmpty;
  wire T32;
  wire T33;
  wire T34;
  wire[31:0] T35;
  reg [31:0] ram [1:0];
  wire[31:0] T36;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    isFull = {1{$random}};
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_enqRdyOut = T0;
  assign T0 = T1 & io_enqValid;
  assign T1 = isFull ^ 1'h1;
  assign T37 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T4 ? 1'h1 : T2;
  assign T2 = T3 ? 1'h0 : isFull;
  assign T3 = doDeq & isFull;
  assign doDeq = io_deqValid;
  assign T4 = T10 & T5;
  assign T5 = enqPtrInc == deqPtr;
  assign T38 = reset ? 1'h0 : T6;
  assign T6 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T7 % 2'h2;
  assign T7 = deqPtr + 1'h1;
  assign enqPtrInc = T8 % 2'h2;
  assign T8 = enqPtr + 1'h1;
  assign T39 = reset ? 1'h0 : T9;
  assign T9 = doEnq ? enqPtrInc : enqPtr;
  assign doEnq = io_enqRdyOut;
  assign T10 = doEnq & T11;
  assign T11 = ~ doDeq;
  assign io_deqValid = T12;
  assign T12 = T31 & deqCombined;
  assign deqCombined = deqCond == 4'hf;
  assign deqCond = {T22, T13};
  assign T13 = {T18, T14};
  assign T14 = T17 | T15;
  assign T15 = ~ T16;
  assign T16 = io_deqReg[2'h3:2'h3];
  assign T17 = io_deqRdy[2'h3:2'h3];
  assign T18 = T21 | T19;
  assign T19 = ~ T20;
  assign T20 = io_deqReg[2'h2:2'h2];
  assign T21 = io_deqRdy[2'h2:2'h2];
  assign T22 = {T27, T23};
  assign T23 = T26 | T24;
  assign T24 = ~ T25;
  assign T25 = io_deqReg[1'h1:1'h1];
  assign T26 = io_deqRdy[1'h1:1'h1];
  assign T27 = T30 | T28;
  assign T28 = ~ T29;
  assign T29 = io_deqReg[1'h0:1'h0];
  assign T30 = io_deqRdy[1'h0:1'h0];
  assign T31 = isEmpty ^ 1'h1;
  assign isEmpty = T33 & T32;
  assign T32 = enqPtr == deqPtr;
  assign T33 = isFull ^ 1'h1;
  assign io_enqRdy = T34;
  assign T34 = isFull ^ 1'h1;
  assign io_deqData = T35;
  assign T35 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      isFull <= 1'h0;
    end else if(T4) begin
      isFull <= 1'h1;
    end else if(T3) begin
      isFull <= 1'h0;
    end
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Mux_0(
    input [32:0] io_inMuxPort_3,
    input [32:0] io_inMuxPort_2,
    input [32:0] io_inMuxPort_1,
    input [32:0] io_inMuxPort_0,
    input [1:0] io_sel,
    output[31:0] io_outMuxPort
);

  wire[31:0] T7;
  wire[32:0] T0;
  wire[32:0] T1;
  wire T2;
  wire[1:0] T3;
  wire[32:0] T4;
  wire T5;
  wire T6;


  assign io_outMuxPort = T7;
  assign T7 = T0[5'h1f:1'h0];
  assign T0 = T6 ? T4 : T1;
  assign T1 = T2 ? io_inMuxPort_1 : io_inMuxPort_0;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = io_sel;
  assign T4 = T5 ? io_inMuxPort_3 : io_inMuxPort_2;
  assign T5 = T3[1'h0:1'h0];
  assign T6 = T3[1'h1:1'h1];
endmodule

module Mux_1(
    input  io_inMuxPort_3,
    input  io_inMuxPort_2,
    input  io_inMuxPort_1,
    input  io_inMuxPort_0,
    input [1:0] io_sel,
    output io_outMuxPort
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_outMuxPort = T0;
  assign T0 = T6 ? T4 : T1;
  assign T1 = T2 ? io_inMuxPort_1 : io_inMuxPort_0;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = io_sel;
  assign T4 = T5 ? io_inMuxPort_3 : io_inMuxPort_2;
  assign T5 = T3[1'h0:1'h0];
  assign T6 = T3[1'h1:1'h1];
endmodule

module CU(input clk, input reset,
    input [32:0] io_in_3,
    input [32:0] io_in_2,
    input [32:0] io_in_1,
    input [32:0] io_in_0,
    output[32:0] io_out,
    input [23:0] io_inConfig,
    output io_enqRdy,
    input [3:0] io_deqRdy,
    input [3:0] io_enqValid,
    output io_deqValid,
    output io_enqRdyOut
);

  wire[1:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire[31:0] T23;
  wire[32:0] T15;
  wire[32:0] T16;
  wire T17;
  wire T18;
  wire[4:0] T24;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[32:0] T25;
  wire[31:0] ALUClass_io_out;
  wire ALUClass_io_outValid;
  wire[31:0] FifoCUClass_io_deqData;
  wire FifoCUClass_io_enqRdy;
  wire FifoCUClass_io_deqValid;
  wire FifoCUClass_io_enqRdyOut;
  wire[31:0] MuxIn1_io_outMuxPort;
  wire[31:0] MuxIn2_io_outMuxPort;
  wire MuxInValid1_io_outMuxPort;
  wire MuxInValid2_io_outMuxPort;


  assign T0 = io_inConfig[4'h8:3'h7];
  assign T1 = io_enqValid[1'h0:1'h0];
  assign T2 = io_enqValid[1'h1:1'h1];
  assign T3 = io_enqValid[2'h2:2'h2];
  assign T4 = io_enqValid[2'h3:2'h3];
  assign T5 = io_inConfig[3'h6:3'h5];
  assign T6 = io_enqValid[1'h0:1'h0];
  assign T7 = io_enqValid[1'h1:1'h1];
  assign T8 = io_enqValid[2'h2:2'h2];
  assign T9 = io_enqValid[2'h3:2'h3];
  assign T10 = io_inConfig[4'h8:3'h7];
  assign T11 = io_inConfig[3'h6:3'h5];
  assign T12 = io_inConfig[4'hc:4'h9];
  assign T13 = T14 ? 1'h0 : ALUClass_io_outValid;
  assign T14 = io_inConfig[3'h4:3'h4];
  assign T23 = T15[5'h1f:1'h0];
  assign T15 = T14 ? 33'h0 : T16;
  assign T16 = {1'h0, ALUClass_io_out};
  assign T17 = T14 ? 1'h0 : MuxInValid2_io_outMuxPort;
  assign T18 = T14 ? 1'h0 : MuxInValid1_io_outMuxPort;
  assign T24 = {1'h0, T19};
  assign T19 = T14 ? 4'hf : T20;
  assign T20 = io_inConfig[2'h3:1'h0];
  assign T21 = T14 ? 32'h0 : MuxIn2_io_outMuxPort;
  assign T22 = T14 ? 32'h0 : MuxIn1_io_outMuxPort;
  assign io_enqRdyOut = FifoCUClass_io_enqRdyOut;
  assign io_deqValid = FifoCUClass_io_deqValid;
  assign io_enqRdy = FifoCUClass_io_enqRdy;
  assign io_out = T25;
  assign T25 = {1'h0, FifoCUClass_io_deqData};
  ALU ALUClass(
       .io_inOp1( T22 ),
       .io_inOp2( T21 ),
       .io_out( ALUClass_io_out ),
       .io_opCode( T24 ),
       .io_inOp1Valid( T18 ),
       .io_inOp2Valid( T17 ),
       .io_outValid( ALUClass_io_outValid )
  );
  FifoCU FifoCUClass(.clk(clk), .reset(reset),
       .io_enqData( T23 ),
       .io_deqData( FifoCUClass_io_deqData ),
       .io_enqRdy( FifoCUClass_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( T13 ),
       .io_deqValid( FifoCUClass_io_deqValid ),
       .io_deqReg( T12 ),
       .io_enqRdyOut( FifoCUClass_io_enqRdyOut )
  );
  Mux_0 MuxIn1(
       .io_inMuxPort_3( io_in_3 ),
       .io_inMuxPort_2( io_in_2 ),
       .io_inMuxPort_1( io_in_1 ),
       .io_inMuxPort_0( io_in_0 ),
       .io_sel( T11 ),
       .io_outMuxPort( MuxIn1_io_outMuxPort )
  );
  Mux_0 MuxIn2(
       .io_inMuxPort_3( io_in_3 ),
       .io_inMuxPort_2( io_in_2 ),
       .io_inMuxPort_1( io_in_1 ),
       .io_inMuxPort_0( io_in_0 ),
       .io_sel( T10 ),
       .io_outMuxPort( MuxIn2_io_outMuxPort )
  );
  Mux_1 MuxInValid1(
       .io_inMuxPort_3( T9 ),
       .io_inMuxPort_2( T8 ),
       .io_inMuxPort_1( T7 ),
       .io_inMuxPort_0( T6 ),
       .io_sel( T5 ),
       .io_outMuxPort( MuxInValid1_io_outMuxPort )
  );
  Mux_1 MuxInValid2(
       .io_inMuxPort_3( T4 ),
       .io_inMuxPort_2( T3 ),
       .io_inMuxPort_1( T2 ),
       .io_inMuxPort_0( T1 ),
       .io_sel( T0 ),
       .io_outMuxPort( MuxInValid2_io_outMuxPort )
  );
endmodule

module Fifo_0(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h0;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_1(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h1;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_2(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h2;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_3(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h3;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_4(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h4;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_5(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h5;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_6(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h6;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module Fifo_7(input clk, input reset,
    input [32:0] io_enqData,
    output[32:0] io_deqData,
    output io_enqRdy,
    input [7:0] io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input [23:0] io_configVal,
    input  io_deqOR
);

  wire T0;
  wire deqCombined;
  wire T1;
  wire[7:0] deqCond;
  wire[3:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire deqReg_7;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] ownReg;
  wire T13;
  wire T14;
  wire T15;
  wire deqReg_6;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire deqReg_5;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire deqReg_4;
  wire T37;
  wire T38;
  wire[2:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire deqReg_3;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire deqReg_2;
  wire T59;
  wire T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire deqReg_1;
  wire T70;
  wire T71;
  wire[2:0] T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire deqReg_0;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire isEmpty;
  wire T90;
  reg  deqPtr;
  wire T106;
  wire T91;
  wire deqPtrInc;
  wire T92;
  wire doDeq;
  reg  enqPtr;
  wire T107;
  wire T93;
  wire enqPtrInc;
  wire T94;
  wire doEnq;
  wire T95;
  wire T96;
  reg  isFull;
  wire T108;
  wire isFullNext;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[32:0] T104;
  reg [32:0] ram [1:0];
  wire[32:0] T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = T89 & deqCombined;
  assign deqCombined = io_deqOR ? T88 : T1;
  assign T1 = deqCond == 8'hff;
  assign deqCond = {T45, T2};
  assign T2 = {T24, T3};
  assign T3 = {T14, T4};
  assign T4 = T13 | T5;
  assign T5 = ~ deqReg_7;
  assign deqReg_7 = T6;
  assign T6 = T7 ? 1'h1 : 1'h0;
  assign T7 = ownReg == T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = io_configVal[5'h15:5'h15];
  assign T11 = io_configVal[5'h16:5'h16];
  assign T12 = io_configVal[5'h17:5'h17];
  assign ownReg = 3'h7;
  assign T13 = io_deqRdy[3'h7:3'h7];
  assign T14 = T23 | T15;
  assign T15 = ~ deqReg_6;
  assign deqReg_6 = T16;
  assign T16 = T17 ? 1'h1 : 1'h0;
  assign T17 = ownReg == T18;
  assign T18 = {T22, T19};
  assign T19 = {T21, T20};
  assign T20 = io_configVal[5'h12:5'h12];
  assign T21 = io_configVal[5'h13:5'h13];
  assign T22 = io_configVal[5'h14:5'h14];
  assign T23 = io_deqRdy[3'h6:3'h6];
  assign T24 = {T35, T25};
  assign T25 = T34 | T26;
  assign T26 = ~ deqReg_5;
  assign deqReg_5 = T27;
  assign T27 = T28 ? 1'h1 : 1'h0;
  assign T28 = ownReg == T29;
  assign T29 = {T33, T30};
  assign T30 = {T32, T31};
  assign T31 = io_configVal[4'hf:4'hf];
  assign T32 = io_configVal[5'h10:5'h10];
  assign T33 = io_configVal[5'h11:5'h11];
  assign T34 = io_deqRdy[3'h5:3'h5];
  assign T35 = T44 | T36;
  assign T36 = ~ deqReg_4;
  assign deqReg_4 = T37;
  assign T37 = T38 ? 1'h1 : 1'h0;
  assign T38 = ownReg == T39;
  assign T39 = {T43, T40};
  assign T40 = {T42, T41};
  assign T41 = io_configVal[4'hc:4'hc];
  assign T42 = io_configVal[4'hd:4'hd];
  assign T43 = io_configVal[4'he:4'he];
  assign T44 = io_deqRdy[3'h4:3'h4];
  assign T45 = {T67, T46};
  assign T46 = {T57, T47};
  assign T47 = T56 | T48;
  assign T48 = ~ deqReg_3;
  assign deqReg_3 = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = ownReg == T51;
  assign T51 = {T55, T52};
  assign T52 = {T54, T53};
  assign T53 = io_configVal[4'h9:4'h9];
  assign T54 = io_configVal[4'ha:4'ha];
  assign T55 = io_configVal[4'hb:4'hb];
  assign T56 = io_deqRdy[2'h3:2'h3];
  assign T57 = T66 | T58;
  assign T58 = ~ deqReg_2;
  assign deqReg_2 = T59;
  assign T59 = T60 ? 1'h1 : 1'h0;
  assign T60 = ownReg == T61;
  assign T61 = {T65, T62};
  assign T62 = {T64, T63};
  assign T63 = io_configVal[3'h6:3'h6];
  assign T64 = io_configVal[3'h7:3'h7];
  assign T65 = io_configVal[4'h8:4'h8];
  assign T66 = io_deqRdy[2'h2:2'h2];
  assign T67 = {T78, T68};
  assign T68 = T77 | T69;
  assign T69 = ~ deqReg_1;
  assign deqReg_1 = T70;
  assign T70 = T71 ? 1'h1 : 1'h0;
  assign T71 = ownReg == T72;
  assign T72 = {T76, T73};
  assign T73 = {T75, T74};
  assign T74 = io_configVal[2'h3:2'h3];
  assign T75 = io_configVal[3'h4:3'h4];
  assign T76 = io_configVal[3'h5:3'h5];
  assign T77 = io_deqRdy[1'h1:1'h1];
  assign T78 = T87 | T79;
  assign T79 = ~ deqReg_0;
  assign deqReg_0 = T80;
  assign T80 = T81 ? 1'h1 : 1'h0;
  assign T81 = ownReg == T82;
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = io_configVal[1'h0:1'h0];
  assign T85 = io_configVal[1'h1:1'h1];
  assign T86 = io_configVal[2'h2:2'h2];
  assign T87 = io_deqRdy[1'h0:1'h0];
  assign T88 = io_deqRdy[1'h1:1'h1];
  assign T89 = isEmpty ^ 1'h1;
  assign isEmpty = T96 & T90;
  assign T90 = enqPtr == deqPtr;
  assign T106 = reset ? 1'h0 : T91;
  assign T91 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T92 % 2'h2;
  assign T92 = deqPtr + 1'h1;
  assign doDeq = io_deqValid;
  assign T107 = reset ? 1'h0 : T93;
  assign T93 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T94 % 2'h2;
  assign T94 = enqPtr + 1'h1;
  assign doEnq = T95;
  assign T95 = io_enqRdy & io_enqValid;
  assign T96 = isFull ^ 1'h1;
  assign T108 = reset ? 1'h0 : isFullNext;
  assign isFullNext = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : isFull;
  assign T98 = doDeq & isFull;
  assign T99 = T101 & T100;
  assign T100 = enqPtrInc == deqPtr;
  assign T101 = doEnq & T102;
  assign T102 = ~ doDeq;
  assign io_enqRdy = T103;
  assign T103 = isFull ^ 1'h1;
  assign io_deqData = T104;
  assign T104 = ram[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(T99) begin
      isFull <= 1'h1;
    end else if(T98) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      ram[enqPtr] <= io_enqData;
  end
endmodule

module MuxSwitch_0(
    input [32:0] io_inMuxPort_7,
    input [32:0] io_inMuxPort_6,
    input [32:0] io_inMuxPort_5,
    input [32:0] io_inMuxPort_4,
    input [32:0] io_inMuxPort_3,
    input [32:0] io_inMuxPort_2,
    input [32:0] io_inMuxPort_1,
    input [32:0] io_inMuxPort_0,
    input [2:0] io_sel,
    output[32:0] io_outMuxPort
);

  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[32:0] T5;
  wire T6;
  wire T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire T10;
  wire[32:0] T11;
  wire T12;
  wire T13;
  wire T14;


  assign io_outMuxPort = T0;
  assign T0 = T14 ? T8 : T1;
  assign T1 = T7 ? T5 : T2;
  assign T2 = T3 ? io_inMuxPort_1 : io_inMuxPort_0;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = io_sel;
  assign T5 = T6 ? io_inMuxPort_3 : io_inMuxPort_2;
  assign T6 = T4[1'h0:1'h0];
  assign T7 = T4[1'h1:1'h1];
  assign T8 = T13 ? T11 : T9;
  assign T9 = T10 ? io_inMuxPort_5 : io_inMuxPort_4;
  assign T10 = T4[1'h0:1'h0];
  assign T11 = T12 ? io_inMuxPort_7 : io_inMuxPort_6;
  assign T12 = T4[1'h0:1'h0];
  assign T13 = T4[1'h1:1'h1];
  assign T14 = T4[2'h2:2'h2];
endmodule

module MuxSwitch_1(
    input  io_inMuxPort_7,
    input  io_inMuxPort_6,
    input  io_inMuxPort_5,
    input  io_inMuxPort_4,
    input  io_inMuxPort_3,
    input  io_inMuxPort_2,
    input  io_inMuxPort_1,
    input  io_inMuxPort_0,
    input [2:0] io_sel,
    output io_outMuxPort
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;


  assign io_outMuxPort = T0;
  assign T0 = T14 ? T8 : T1;
  assign T1 = T7 ? T5 : T2;
  assign T2 = T3 ? io_inMuxPort_1 : io_inMuxPort_0;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = io_sel;
  assign T5 = T6 ? io_inMuxPort_3 : io_inMuxPort_2;
  assign T6 = T4[1'h0:1'h0];
  assign T7 = T4[1'h1:1'h1];
  assign T8 = T13 ? T11 : T9;
  assign T9 = T10 ? io_inMuxPort_5 : io_inMuxPort_4;
  assign T10 = T4[1'h0:1'h0];
  assign T11 = T12 ? io_inMuxPort_7 : io_inMuxPort_6;
  assign T12 = T4[1'h0:1'h0];
  assign T13 = T4[1'h1:1'h1];
  assign T14 = T4[2'h2:2'h2];
endmodule

module Crossbar(
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    input [23:0] io_inSwitchConfig,
    input  io_enqValidIn_7,
    input  io_enqValidIn_6,
    input  io_enqValidIn_5,
    input  io_enqValidIn_4,
    input  io_enqValidIn_3,
    input  io_enqValidIn_2,
    input  io_enqValidIn_1,
    input  io_enqValidIn_0,
    output io_enqValidOut_7,
    output io_enqValidOut_6,
    output io_enqValidOut_5,
    output io_enqValidOut_4,
    output io_enqValidOut_3,
    output io_enqValidOut_2,
    output io_enqValidOut_1,
    output io_enqValidOut_0,
    input [32:0] io_inConfigData,
    input  io_enqConfigPort_1
);

  wire[2:0] T0;
  wire[1:0] T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire[2:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire[2:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire[2:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire[2:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire[2:0] T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[2:0] T65;
  wire[1:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[2:0] T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire[1:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[32:0] T81;
  wire[32:0] MuxSwitch_io_outMuxPort;
  wire[32:0] MuxSwitch_1_io_outMuxPort;
  wire[32:0] MuxSwitch_2_io_outMuxPort;
  wire[32:0] MuxSwitch_3_io_outMuxPort;
  wire[32:0] MuxSwitch_4_io_outMuxPort;
  wire[32:0] MuxSwitch_5_io_outMuxPort;
  wire[32:0] MuxSwitch_6_io_outMuxPort;
  wire[32:0] MuxSwitch_7_io_outMuxPort;
  wire MuxSwitch_8_io_outMuxPort;
  wire MuxSwitch_9_io_outMuxPort;
  wire MuxSwitch_10_io_outMuxPort;
  wire MuxSwitch_11_io_outMuxPort;
  wire MuxSwitch_12_io_outMuxPort;
  wire MuxSwitch_13_io_outMuxPort;
  wire MuxSwitch_14_io_outMuxPort;
  wire MuxSwitch_15_io_outMuxPort;


  assign T0 = {T4, T1};
  assign T1 = {T3, T2};
  assign T2 = io_inSwitchConfig[5'h15:5'h15];
  assign T3 = io_inSwitchConfig[5'h16:5'h16];
  assign T4 = io_inSwitchConfig[5'h17:5'h17];
  assign T5 = {T9, T6};
  assign T6 = {T8, T7};
  assign T7 = io_inSwitchConfig[5'h12:5'h12];
  assign T8 = io_inSwitchConfig[5'h13:5'h13];
  assign T9 = io_inSwitchConfig[5'h14:5'h14];
  assign T10 = {T14, T11};
  assign T11 = {T13, T12};
  assign T12 = io_inSwitchConfig[4'hf:4'hf];
  assign T13 = io_inSwitchConfig[5'h10:5'h10];
  assign T14 = io_inSwitchConfig[5'h11:5'h11];
  assign T15 = {T19, T16};
  assign T16 = {T18, T17};
  assign T17 = io_inSwitchConfig[4'hc:4'hc];
  assign T18 = io_inSwitchConfig[4'hd:4'hd];
  assign T19 = io_inSwitchConfig[4'he:4'he];
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_inSwitchConfig[4'h9:4'h9];
  assign T23 = io_inSwitchConfig[4'ha:4'ha];
  assign T24 = io_inSwitchConfig[4'hb:4'hb];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_inSwitchConfig[3'h6:3'h6];
  assign T28 = io_inSwitchConfig[3'h7:3'h7];
  assign T29 = io_inSwitchConfig[4'h8:4'h8];
  assign T30 = {T34, T31};
  assign T31 = {T33, T32};
  assign T32 = io_inSwitchConfig[2'h3:2'h3];
  assign T33 = io_inSwitchConfig[3'h4:3'h4];
  assign T34 = io_inSwitchConfig[3'h5:3'h5];
  assign T35 = {T39, T36};
  assign T36 = {T38, T37};
  assign T37 = io_inSwitchConfig[1'h0:1'h0];
  assign T38 = io_inSwitchConfig[1'h1:1'h1];
  assign T39 = io_inSwitchConfig[2'h2:2'h2];
  assign T40 = {T44, T41};
  assign T41 = {T43, T42};
  assign T42 = io_inSwitchConfig[5'h15:5'h15];
  assign T43 = io_inSwitchConfig[5'h16:5'h16];
  assign T44 = io_inSwitchConfig[5'h17:5'h17];
  assign T45 = {T49, T46};
  assign T46 = {T48, T47};
  assign T47 = io_inSwitchConfig[5'h12:5'h12];
  assign T48 = io_inSwitchConfig[5'h13:5'h13];
  assign T49 = io_inSwitchConfig[5'h14:5'h14];
  assign T50 = {T54, T51};
  assign T51 = {T53, T52};
  assign T52 = io_inSwitchConfig[4'hf:4'hf];
  assign T53 = io_inSwitchConfig[5'h10:5'h10];
  assign T54 = io_inSwitchConfig[5'h11:5'h11];
  assign T55 = {T59, T56};
  assign T56 = {T58, T57};
  assign T57 = io_inSwitchConfig[4'hc:4'hc];
  assign T58 = io_inSwitchConfig[4'hd:4'hd];
  assign T59 = io_inSwitchConfig[4'he:4'he];
  assign T60 = {T64, T61};
  assign T61 = {T63, T62};
  assign T62 = io_inSwitchConfig[4'h9:4'h9];
  assign T63 = io_inSwitchConfig[4'ha:4'ha];
  assign T64 = io_inSwitchConfig[4'hb:4'hb];
  assign T65 = {T69, T66};
  assign T66 = {T68, T67};
  assign T67 = io_inSwitchConfig[3'h6:3'h6];
  assign T68 = io_inSwitchConfig[3'h7:3'h7];
  assign T69 = io_inSwitchConfig[4'h8:4'h8];
  assign T70 = {T74, T71};
  assign T71 = {T73, T72};
  assign T72 = io_inSwitchConfig[2'h3:2'h3];
  assign T73 = io_inSwitchConfig[3'h4:3'h4];
  assign T74 = io_inSwitchConfig[3'h5:3'h5];
  assign T75 = {T79, T76};
  assign T76 = {T78, T77};
  assign T77 = io_inSwitchConfig[1'h0:1'h0];
  assign T78 = io_inSwitchConfig[1'h1:1'h1];
  assign T79 = io_inSwitchConfig[2'h2:2'h2];
  assign io_enqValidOut_0 = MuxSwitch_8_io_outMuxPort;
  assign io_enqValidOut_1 = T80;
  assign T80 = io_enqConfigPort_1 ? io_enqConfigPort_1 : MuxSwitch_9_io_outMuxPort;
  assign io_enqValidOut_2 = MuxSwitch_10_io_outMuxPort;
  assign io_enqValidOut_3 = MuxSwitch_11_io_outMuxPort;
  assign io_enqValidOut_4 = MuxSwitch_12_io_outMuxPort;
  assign io_enqValidOut_5 = MuxSwitch_13_io_outMuxPort;
  assign io_enqValidOut_6 = MuxSwitch_14_io_outMuxPort;
  assign io_enqValidOut_7 = MuxSwitch_15_io_outMuxPort;
  assign io_outPort_0 = MuxSwitch_io_outMuxPort;
  assign io_outPort_1 = T81;
  assign T81 = io_enqConfigPort_1 ? io_inConfigData : MuxSwitch_1_io_outMuxPort;
  assign io_outPort_2 = MuxSwitch_2_io_outMuxPort;
  assign io_outPort_3 = MuxSwitch_3_io_outMuxPort;
  assign io_outPort_4 = MuxSwitch_4_io_outMuxPort;
  assign io_outPort_5 = MuxSwitch_5_io_outMuxPort;
  assign io_outPort_6 = MuxSwitch_6_io_outMuxPort;
  assign io_outPort_7 = MuxSwitch_7_io_outMuxPort;
  MuxSwitch_0 MuxSwitch(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       //.io_inMuxPort_0(  )
       .io_sel( T75 ),
       .io_outMuxPort( MuxSwitch_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch.io_inMuxPort_0 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_1(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       //.io_inMuxPort_1(  )
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T70 ),
       .io_outMuxPort( MuxSwitch_1_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_1.io_inMuxPort_1 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_2(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       //.io_inMuxPort_2(  )
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T65 ),
       .io_outMuxPort( MuxSwitch_2_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_2.io_inMuxPort_2 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_3(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       //.io_inMuxPort_3(  )
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T60 ),
       .io_outMuxPort( MuxSwitch_3_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_3.io_inMuxPort_3 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_4(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       //.io_inMuxPort_4(  )
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T55 ),
       .io_outMuxPort( MuxSwitch_4_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_4.io_inMuxPort_4 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_5(
       .io_inMuxPort_7( io_inPort_7 ),
       .io_inMuxPort_6( io_inPort_6 ),
       //.io_inMuxPort_5(  )
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T50 ),
       .io_outMuxPort( MuxSwitch_5_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_5.io_inMuxPort_5 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_6(
       .io_inMuxPort_7( io_inPort_7 ),
       //.io_inMuxPort_6(  )
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T45 ),
       .io_outMuxPort( MuxSwitch_6_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_6.io_inMuxPort_6 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_0 MuxSwitch_7(
       //.io_inMuxPort_7(  )
       .io_inMuxPort_6( io_inPort_6 ),
       .io_inMuxPort_5( io_inPort_5 ),
       .io_inMuxPort_4( io_inPort_4 ),
       .io_inMuxPort_3( io_inPort_3 ),
       .io_inMuxPort_2( io_inPort_2 ),
       .io_inMuxPort_1( io_inPort_1 ),
       .io_inMuxPort_0( io_inPort_0 ),
       .io_sel( T40 ),
       .io_outMuxPort( MuxSwitch_7_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_7.io_inMuxPort_7 = {2{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_8(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       //.io_inMuxPort_0(  )
       .io_sel( T35 ),
       .io_outMuxPort( MuxSwitch_8_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_8.io_inMuxPort_0 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_9(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       //.io_inMuxPort_1(  )
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T30 ),
       .io_outMuxPort( MuxSwitch_9_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_9.io_inMuxPort_1 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_10(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       //.io_inMuxPort_2(  )
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T25 ),
       .io_outMuxPort( MuxSwitch_10_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_10.io_inMuxPort_2 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_11(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       //.io_inMuxPort_3(  )
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T20 ),
       .io_outMuxPort( MuxSwitch_11_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_11.io_inMuxPort_3 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_12(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       //.io_inMuxPort_4(  )
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T15 ),
       .io_outMuxPort( MuxSwitch_12_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_12.io_inMuxPort_4 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_13(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       .io_inMuxPort_6( io_enqValidIn_6 ),
       //.io_inMuxPort_5(  )
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T10 ),
       .io_outMuxPort( MuxSwitch_13_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_13.io_inMuxPort_5 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_14(
       .io_inMuxPort_7( io_enqValidIn_7 ),
       //.io_inMuxPort_6(  )
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T5 ),
       .io_outMuxPort( MuxSwitch_14_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_14.io_inMuxPort_6 = {1{$random}};
// synthesis translate_on
`endif
  MuxSwitch_1 MuxSwitch_15(
       //.io_inMuxPort_7(  )
       .io_inMuxPort_6( io_enqValidIn_6 ),
       .io_inMuxPort_5( io_enqValidIn_5 ),
       .io_inMuxPort_4( io_enqValidIn_4 ),
       .io_inMuxPort_3( io_enqValidIn_3 ),
       .io_inMuxPort_2( io_enqValidIn_2 ),
       .io_inMuxPort_1( io_enqValidIn_1 ),
       .io_inMuxPort_0( io_enqValidIn_0 ),
       .io_sel( T0 ),
       .io_outMuxPort( MuxSwitch_15_io_outMuxPort )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxSwitch_15.io_inMuxPort_7 = {1{$random}};
// synthesis translate_on
`endif
endmodule

module Switch_0(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h0;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module Switch_1(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h1;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module Switch_2(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h2;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module Switch_3(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h3;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module Switch_4(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h4;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module Switch_5(input clk, input reset,
    input [32:0] io_inPort_7,
    input [32:0] io_inPort_6,
    input [32:0] io_inPort_5,
    input [32:0] io_inPort_4,
    input [32:0] io_inPort_3,
    input [32:0] io_inPort_2,
    input [32:0] io_inPort_1,
    input [32:0] io_inPort_0,
    output[32:0] io_outPort_7,
    output[32:0] io_outPort_6,
    output[32:0] io_outPort_5,
    output[32:0] io_outPort_4,
    output[32:0] io_outPort_3,
    output[32:0] io_outPort_2,
    output[32:0] io_outPort_1,
    output[32:0] io_outPort_0,
    output[7:0] io_deqValid,
    output[7:0] io_enqRdy,
    input [7:0] io_deqRdy,
    input [7:0] io_enqValid,
    output[32:0] io_outConfigData,
    output[23:0] io_outCUConfig,
    input  io_deqOR,
    output io_enqOR,
    input [3:0] io_deqRdyOut
);

  wire enqConfigPort_1;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] inYCoord;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire T7;
  wire[32:0] inConfigData;
  wire[32:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire inType;
  wire T12;
  wire[32:0] inCheckData;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[7:0] enqValidTweaked;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg [23:0] sConfigReg;
  wire[23:0] T178;
  wire[23:0] T39;
  wire[23:0] T40;
  wire[11:0] T41;
  wire[5:0] T42;
  wire[2:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[5:0] T53;
  wire[2:0] T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire[11:0] T64;
  wire[5:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[2:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[5:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire configType;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[6:0] T93;
  wire T94;
  wire[7:0] T95;
  wire[6:0] T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire[7:0] T100;
  wire[5:0] T101;
  wire[4:0] T102;
  wire T103;
  wire[1:0] T104;
  wire[7:0] T105;
  wire[4:0] T106;
  wire[3:0] T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  reg [23:0] cuConfigReg;
  wire[23:0] T179;
  wire[23:0] T114;
  wire[23:0] T115;
  wire[11:0] T116;
  wire[5:0] T117;
  wire[2:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire[2:0] T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[5:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[11:0] T139;
  wire[5:0] T140;
  wire[2:0] T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[2:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire T150;
  wire[5:0] T151;
  wire[2:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[2:0] T157;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[7:0] T171;
  wire[3:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[3:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[32:0] Fifo_io_deqData;
  wire Fifo_io_enqRdy;
  wire Fifo_io_deqValid;
  wire[32:0] Fifo_1_io_deqData;
  wire Fifo_1_io_enqRdy;
  wire Fifo_1_io_deqValid;
  wire[32:0] Fifo_2_io_deqData;
  wire Fifo_2_io_enqRdy;
  wire Fifo_2_io_deqValid;
  wire[32:0] Fifo_3_io_deqData;
  wire Fifo_3_io_enqRdy;
  wire Fifo_3_io_deqValid;
  wire[32:0] Fifo_4_io_deqData;
  wire Fifo_4_io_enqRdy;
  wire Fifo_4_io_deqValid;
  wire[32:0] Fifo_5_io_deqData;
  wire Fifo_5_io_enqRdy;
  wire Fifo_5_io_deqValid;
  wire[32:0] Fifo_6_io_deqData;
  wire Fifo_6_io_enqRdy;
  wire Fifo_6_io_deqValid;
  wire[32:0] Fifo_7_io_deqData;
  wire Fifo_7_io_enqRdy;
  wire Fifo_7_io_deqValid;
  wire[32:0] crossbarClass_io_outPort_7;
  wire[32:0] crossbarClass_io_outPort_6;
  wire[32:0] crossbarClass_io_outPort_5;
  wire[32:0] crossbarClass_io_outPort_4;
  wire[32:0] crossbarClass_io_outPort_3;
  wire[32:0] crossbarClass_io_outPort_2;
  wire[32:0] crossbarClass_io_outPort_1;
  wire[32:0] crossbarClass_io_outPort_0;
  wire crossbarClass_io_enqValidOut_7;
  wire crossbarClass_io_enqValidOut_6;
  wire crossbarClass_io_enqValidOut_5;
  wire crossbarClass_io_enqValidOut_4;
  wire crossbarClass_io_enqValidOut_3;
  wire crossbarClass_io_enqValidOut_2;
  wire crossbarClass_io_enqValidOut_1;
  wire crossbarClass_io_enqValidOut_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sConfigReg = {1{$random}};
    cuConfigReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign enqConfigPort_1 = T0;
  assign T0 = T14 ? T13 : T1;
  assign T1 = T2 ? 1'h0 : 1'h0;
  assign T2 = T11 & T3;
  assign T3 = inYCoord == 3'h5;
  assign inYCoord = T4;
  assign T4 = T11 ? T5 : 3'h0;
  assign T5 = {T10, T6};
  assign T6 = {T9, T7};
  assign T7 = inConfigData[5'h1d:5'h1d];
  assign inConfigData = T8;
  assign T8 = T11 ? io_inPort_3 : 33'h0;
  assign T9 = inConfigData[5'h1e:5'h1e];
  assign T10 = inConfigData[5'h1f:5'h1f];
  assign T11 = inType;
  assign inType = T12;
  assign T12 = inCheckData[6'h20:6'h20];
  assign inCheckData = io_inPort_3;
  assign T13 = io_enqValid[2'h3:2'h3];
  assign T14 = T11 & T15;
  assign T15 = T3 ^ 1'h1;
  assign T16 = enqValidTweaked[1'h0:1'h0];
  assign enqValidTweaked = T17;
  assign T17 = T11 ? T18 : io_enqValid;
  assign T18 = {T25, T19};
  assign T19 = {1'h0, T20};
  assign T20 = {T24, T21};
  assign T21 = {T23, T22};
  assign T22 = io_enqValid[1'h0:1'h0];
  assign T23 = io_enqValid[1'h1:1'h1];
  assign T24 = io_enqValid[2'h2:2'h2];
  assign T25 = {T29, T26};
  assign T26 = {T28, T27};
  assign T27 = io_enqValid[3'h4:3'h4];
  assign T28 = io_enqValid[3'h5:3'h5];
  assign T29 = {T31, T30};
  assign T30 = io_enqValid[3'h6:3'h6];
  assign T31 = io_enqValid[3'h7:3'h7];
  assign T32 = enqValidTweaked[1'h1:1'h1];
  assign T33 = enqValidTweaked[2'h2:2'h2];
  assign T34 = enqValidTweaked[2'h3:2'h3];
  assign T35 = enqValidTweaked[3'h4:3'h4];
  assign T36 = enqValidTweaked[3'h5:3'h5];
  assign T37 = enqValidTweaked[3'h6:3'h6];
  assign T38 = enqValidTweaked[3'h7:3'h7];
  assign T178 = reset ? 24'h0 : T39;
  assign T39 = T87 ? T40 : sConfigReg;
  assign T40 = {T64, T41};
  assign T41 = {T53, T42};
  assign T42 = {T48, T43};
  assign T43 = {T47, T44};
  assign T44 = {T46, T45};
  assign T45 = inConfigData[1'h0:1'h0];
  assign T46 = inConfigData[1'h1:1'h1];
  assign T47 = inConfigData[2'h2:2'h2];
  assign T48 = {T52, T49};
  assign T49 = {T51, T50};
  assign T50 = inConfigData[2'h3:2'h3];
  assign T51 = inConfigData[3'h4:3'h4];
  assign T52 = inConfigData[3'h5:3'h5];
  assign T53 = {T59, T54};
  assign T54 = {T58, T55};
  assign T55 = {T57, T56};
  assign T56 = inConfigData[3'h6:3'h6];
  assign T57 = inConfigData[3'h7:3'h7];
  assign T58 = inConfigData[4'h8:4'h8];
  assign T59 = {T63, T60};
  assign T60 = {T62, T61};
  assign T61 = inConfigData[4'h9:4'h9];
  assign T62 = inConfigData[4'ha:4'ha];
  assign T63 = inConfigData[4'hb:4'hb];
  assign T64 = {T76, T65};
  assign T65 = {T71, T66};
  assign T66 = {T70, T67};
  assign T67 = {T69, T68};
  assign T68 = inConfigData[4'hc:4'hc];
  assign T69 = inConfigData[4'hd:4'hd];
  assign T70 = inConfigData[4'he:4'he];
  assign T71 = {T75, T72};
  assign T72 = {T74, T73};
  assign T73 = inConfigData[4'hf:4'hf];
  assign T74 = inConfigData[5'h10:5'h10];
  assign T75 = inConfigData[5'h11:5'h11];
  assign T76 = {T82, T77};
  assign T77 = {T81, T78};
  assign T78 = {T80, T79};
  assign T79 = inConfigData[5'h12:5'h12];
  assign T80 = inConfigData[5'h13:5'h13];
  assign T81 = inConfigData[5'h14:5'h14];
  assign T82 = {T86, T83};
  assign T83 = {T85, T84};
  assign T84 = inConfigData[5'h15:5'h15];
  assign T85 = inConfigData[5'h16:5'h16];
  assign T86 = inConfigData[5'h17:5'h17];
  assign T87 = T2 & T88;
  assign T88 = configType == 1'h1;
  assign configType = T89;
  assign T89 = T14 ? 1'h0 : T90;
  assign T90 = T2 ? T91 : 1'h0;
  assign T91 = inConfigData[5'h1c:5'h1c];
  assign T92 = {T94, T93};
  assign T93 = io_deqRdy[3'h6:1'h0];
  assign T94 = io_deqRdyOut[2'h3:2'h3];
  assign T95 = {T99, T96};
  assign T96 = {T98, T97};
  assign T97 = io_deqRdy[3'h5:1'h0];
  assign T98 = io_deqRdyOut[2'h2:2'h2];
  assign T99 = io_deqRdy[3'h7:3'h7];
  assign T100 = {T104, T101};
  assign T101 = {T103, T102};
  assign T102 = io_deqRdy[3'h4:1'h0];
  assign T103 = io_deqRdyOut[1'h1:1'h1];
  assign T104 = io_deqRdy[3'h7:3'h6];
  assign T105 = {T109, T106};
  assign T106 = {T108, T107};
  assign T107 = io_deqRdy[2'h3:1'h0];
  assign T108 = io_deqRdyOut[1'h0:1'h0];
  assign T109 = io_deqRdy[3'h7:3'h5];
  assign io_enqOR = T110;
  assign T110 = T14 ? T112 : T111;
  assign T111 = T2 ? 1'h1 : 1'h0;
  assign T112 = T113;
  assign T113 = io_enqRdy[1'h1:1'h1];
  assign io_outCUConfig = cuConfigReg;
  assign T179 = reset ? 24'h0 : T114;
  assign T114 = T162 ? T115 : cuConfigReg;
  assign T115 = {T139, T116};
  assign T116 = {T128, T117};
  assign T117 = {T123, T118};
  assign T118 = {T122, T119};
  assign T119 = {T121, T120};
  assign T120 = inConfigData[1'h0:1'h0];
  assign T121 = inConfigData[1'h1:1'h1];
  assign T122 = inConfigData[2'h2:2'h2];
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = inConfigData[2'h3:2'h3];
  assign T126 = inConfigData[3'h4:3'h4];
  assign T127 = inConfigData[3'h5:3'h5];
  assign T128 = {T134, T129};
  assign T129 = {T133, T130};
  assign T130 = {T132, T131};
  assign T131 = inConfigData[3'h6:3'h6];
  assign T132 = inConfigData[3'h7:3'h7];
  assign T133 = inConfigData[4'h8:4'h8];
  assign T134 = {T138, T135};
  assign T135 = {T137, T136};
  assign T136 = inConfigData[4'h9:4'h9];
  assign T137 = inConfigData[4'ha:4'ha];
  assign T138 = inConfigData[4'hb:4'hb];
  assign T139 = {T151, T140};
  assign T140 = {T146, T141};
  assign T141 = {T145, T142};
  assign T142 = {T144, T143};
  assign T143 = inConfigData[4'hc:4'hc];
  assign T144 = inConfigData[4'hd:4'hd];
  assign T145 = inConfigData[4'he:4'he];
  assign T146 = {T150, T147};
  assign T147 = {T149, T148};
  assign T148 = inConfigData[4'hf:4'hf];
  assign T149 = inConfigData[5'h10:5'h10];
  assign T150 = inConfigData[5'h11:5'h11];
  assign T151 = {T157, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = inConfigData[5'h12:5'h12];
  assign T155 = inConfigData[5'h13:5'h13];
  assign T156 = inConfigData[5'h14:5'h14];
  assign T157 = {T161, T158};
  assign T158 = {T160, T159};
  assign T159 = inConfigData[5'h15:5'h15];
  assign T160 = inConfigData[5'h16:5'h16];
  assign T161 = inConfigData[5'h17:5'h17];
  assign T162 = T2 & T163;
  assign T163 = T88 ^ 1'h1;
  assign io_outConfigData = io_inPort_3;
  assign io_enqRdy = T164;
  assign T164 = {T168, T165};
  assign T165 = {T167, T166};
  assign T166 = {Fifo_1_io_enqRdy, Fifo_io_enqRdy};
  assign T167 = {Fifo_3_io_enqRdy, Fifo_2_io_enqRdy};
  assign T168 = {T170, T169};
  assign T169 = {Fifo_5_io_enqRdy, Fifo_4_io_enqRdy};
  assign T170 = {Fifo_7_io_enqRdy, Fifo_6_io_enqRdy};
  assign io_deqValid = T171;
  assign T171 = {T175, T172};
  assign T172 = {T174, T173};
  assign T173 = {Fifo_1_io_deqValid, Fifo_io_deqValid};
  assign T174 = {Fifo_3_io_deqValid, Fifo_2_io_deqValid};
  assign T175 = {T177, T176};
  assign T176 = {Fifo_5_io_deqValid, Fifo_4_io_deqValid};
  assign T177 = {Fifo_7_io_deqValid, Fifo_6_io_deqValid};
  assign io_outPort_0 = Fifo_io_deqData;
  assign io_outPort_1 = Fifo_1_io_deqData;
  assign io_outPort_2 = Fifo_2_io_deqData;
  assign io_outPort_3 = Fifo_3_io_deqData;
  assign io_outPort_4 = Fifo_4_io_deqData;
  assign io_outPort_5 = Fifo_5_io_deqData;
  assign io_outPort_6 = Fifo_6_io_deqData;
  assign io_outPort_7 = Fifo_7_io_deqData;
  Fifo_0 Fifo(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_0 ),
       .io_deqData( Fifo_io_deqData ),
       .io_enqRdy( Fifo_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_0 ),
       .io_deqValid( Fifo_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_1 ),
       .io_deqData( Fifo_1_io_deqData ),
       .io_enqRdy( Fifo_1_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_1 ),
       .io_deqValid( Fifo_1_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( io_deqOR )
  );
  Fifo_2 Fifo_2(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_2 ),
       .io_deqData( Fifo_2_io_deqData ),
       .io_enqRdy( Fifo_2_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_2 ),
       .io_deqValid( Fifo_2_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_3 Fifo_3(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_3 ),
       .io_deqData( Fifo_3_io_deqData ),
       .io_enqRdy( Fifo_3_io_enqRdy ),
       .io_deqRdy( io_deqRdy ),
       .io_enqValid( crossbarClass_io_enqValidOut_3 ),
       .io_deqValid( Fifo_3_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_4 Fifo_4(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_4 ),
       .io_deqData( Fifo_4_io_deqData ),
       .io_enqRdy( Fifo_4_io_enqRdy ),
       .io_deqRdy( T105 ),
       .io_enqValid( crossbarClass_io_enqValidOut_4 ),
       .io_deqValid( Fifo_4_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_5 Fifo_5(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_5 ),
       .io_deqData( Fifo_5_io_deqData ),
       .io_enqRdy( Fifo_5_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( crossbarClass_io_enqValidOut_5 ),
       .io_deqValid( Fifo_5_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_6 Fifo_6(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_6 ),
       .io_deqData( Fifo_6_io_deqData ),
       .io_enqRdy( Fifo_6_io_enqRdy ),
       .io_deqRdy( T95 ),
       .io_enqValid( crossbarClass_io_enqValidOut_6 ),
       .io_deqValid( Fifo_6_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Fifo_7 Fifo_7(.clk(clk), .reset(reset),
       .io_enqData( crossbarClass_io_outPort_7 ),
       .io_deqData( Fifo_7_io_deqData ),
       .io_enqRdy( Fifo_7_io_enqRdy ),
       .io_deqRdy( T92 ),
       .io_enqValid( crossbarClass_io_enqValidOut_7 ),
       .io_deqValid( Fifo_7_io_deqValid ),
       .io_configVal( sConfigReg ),
       .io_deqOR( 1'h0 )
  );
  Crossbar crossbarClass(
       .io_inPort_7( io_inPort_7 ),
       .io_inPort_6( io_inPort_6 ),
       .io_inPort_5( io_inPort_5 ),
       .io_inPort_4( io_inPort_4 ),
       .io_inPort_3( io_inPort_3 ),
       .io_inPort_2( io_inPort_2 ),
       .io_inPort_1( io_inPort_1 ),
       .io_inPort_0( io_inPort_0 ),
       .io_outPort_7( crossbarClass_io_outPort_7 ),
       .io_outPort_6( crossbarClass_io_outPort_6 ),
       .io_outPort_5( crossbarClass_io_outPort_5 ),
       .io_outPort_4( crossbarClass_io_outPort_4 ),
       .io_outPort_3( crossbarClass_io_outPort_3 ),
       .io_outPort_2( crossbarClass_io_outPort_2 ),
       .io_outPort_1( crossbarClass_io_outPort_1 ),
       .io_outPort_0( crossbarClass_io_outPort_0 ),
       .io_inSwitchConfig( sConfigReg ),
       .io_enqValidIn_7( T38 ),
       .io_enqValidIn_6( T37 ),
       .io_enqValidIn_5( T36 ),
       .io_enqValidIn_4( T35 ),
       .io_enqValidIn_3( T34 ),
       .io_enqValidIn_2( T33 ),
       .io_enqValidIn_1( T32 ),
       .io_enqValidIn_0( T16 ),
       .io_enqValidOut_7( crossbarClass_io_enqValidOut_7 ),
       .io_enqValidOut_6( crossbarClass_io_enqValidOut_6 ),
       .io_enqValidOut_5( crossbarClass_io_enqValidOut_5 ),
       .io_enqValidOut_4( crossbarClass_io_enqValidOut_4 ),
       .io_enqValidOut_3( crossbarClass_io_enqValidOut_3 ),
       .io_enqValidOut_2( crossbarClass_io_enqValidOut_2 ),
       .io_enqValidOut_1( crossbarClass_io_enqValidOut_1 ),
       .io_enqValidOut_0( crossbarClass_io_enqValidOut_0 ),
       .io_inConfigData( io_outConfigData ),
       .io_enqConfigPort_1( enqConfigPort_1 )
  );

  always @(posedge clk) begin
    if(reset) begin
      sConfigReg <= 24'h0;
    end else if(T87) begin
      sConfigReg <= T40;
    end
    if(reset) begin
      cuConfigReg <= 24'h0;
    end else if(T162) begin
      cuConfigReg <= T115;
    end
  end
endmodule

module HyperCellFabric(input clk, input reset,
    input [32:0] io_inData_19,
    input [32:0] io_inData_18,
    input [32:0] io_inData_17,
    input [32:0] io_inData_16,
    input [32:0] io_inData_15,
    input [32:0] io_inData_14,
    input [32:0] io_inData_13,
    input [32:0] io_inData_12,
    input [32:0] io_inData_11,
    input [32:0] io_inData_10,
    input [32:0] io_inData_9,
    input [32:0] io_inData_8,
    input [32:0] io_inData_7,
    input [32:0] io_inData_6,
    input [32:0] io_inData_5,
    input [32:0] io_inData_4,
    input [32:0] io_inData_3,
    input [32:0] io_inData_2,
    input [32:0] io_inData_1,
    input [32:0] io_inData_0,
    output[32:0] io_outData_19,
    output[32:0] io_outData_18,
    output[32:0] io_outData_17,
    output[32:0] io_outData_16,
    output[32:0] io_outData_15,
    output[32:0] io_outData_14,
    output[32:0] io_outData_13,
    output[32:0] io_outData_12,
    output[32:0] io_outData_11,
    output[32:0] io_outData_10,
    output[32:0] io_outData_9,
    output[32:0] io_outData_8,
    output[32:0] io_outData_7,
    output[32:0] io_outData_6,
    output[32:0] io_outData_5,
    output[32:0] io_outData_4,
    output[32:0] io_outData_3,
    output[32:0] io_outData_2,
    output[32:0] io_outData_1,
    output[32:0] io_outData_0,
    input  io_enqRdy_19,
    input  io_enqRdy_18,
    input  io_enqRdy_17,
    input  io_enqRdy_16,
    input  io_enqRdy_15,
    input  io_enqRdy_14,
    input  io_enqRdy_13,
    input  io_enqRdy_12,
    input  io_enqRdy_11,
    input  io_enqRdy_10,
    input  io_enqRdy_9,
    input  io_enqRdy_8,
    input  io_enqRdy_7,
    input  io_enqRdy_6,
    input  io_enqRdy_5,
    input  io_enqRdy_4,
    input  io_enqRdy_3,
    input  io_enqRdy_2,
    input  io_enqRdy_1,
    input  io_enqRdy_0,
    input  io_deqValid_19,
    input  io_deqValid_18,
    input  io_deqValid_17,
    input  io_deqValid_16,
    input  io_deqValid_15,
    input  io_deqValid_14,
    input  io_deqValid_13,
    input  io_deqValid_12,
    input  io_deqValid_11,
    input  io_deqValid_10,
    input  io_deqValid_9,
    input  io_deqValid_8,
    input  io_deqValid_7,
    input  io_deqValid_6,
    input  io_deqValid_5,
    input  io_deqValid_4,
    input  io_deqValid_3,
    input  io_deqValid_2,
    input  io_deqValid_1,
    input  io_deqValid_0,
    output io_deqRdy_19,
    output io_deqRdy_18,
    output io_deqRdy_17,
    output io_deqRdy_16,
    output io_deqRdy_15,
    output io_deqRdy_14,
    output io_deqRdy_13,
    output io_deqRdy_12,
    output io_deqRdy_11,
    output io_deqRdy_10,
    output io_deqRdy_9,
    output io_deqRdy_8,
    output io_deqRdy_7,
    output io_deqRdy_6,
    output io_deqRdy_5,
    output io_deqRdy_4,
    output io_deqRdy_3,
    output io_deqRdy_2,
    output io_deqRdy_1,
    output io_deqRdy_0,
    output io_enqValid_19,
    output io_enqValid_18,
    output io_enqValid_17,
    output io_enqValid_16,
    output io_enqValid_15,
    output io_enqValid_14,
    output io_enqValid_13,
    output io_enqValid_12,
    output io_enqValid_11,
    output io_enqValid_10,
    output io_enqValid_9,
    output io_enqValid_8,
    output io_enqValid_7,
    output io_enqValid_6,
    output io_enqValid_5,
    output io_enqValid_4,
    output io_enqValid_3,
    output io_enqValid_2,
    output io_enqValid_1,
    output io_enqValid_0
);

  wire[3:0] T0;
  wire[2:0] T1;
  wire[7:0] T2;
  wire[3:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire[3:0] T8;
  wire[2:0] T9;
  wire[7:0] T10;
  wire[3:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[2:0] T17;
  wire[3:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[7:0] T21;
  wire[3:0] T22;
  wire[1:0] T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[3:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[7:0] T31;
  wire[3:0] T32;
  wire[1:0] T33;
  wire T34;
  wire[1:0] T35;
  wire T36;
  wire T37;
  wire[3:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[3:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[7:0] T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[3:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire[7:0] T54;
  wire[3:0] T55;
  wire[1:0] T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire[3:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire[3:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[7:0] T67;
  wire[3:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire[3:0] T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire[7:0] T77;
  wire[3:0] T78;
  wire[1:0] T79;
  wire T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire[3:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[3:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire[7:0] T90;
  wire[3:0] T91;
  wire[1:0] T92;
  wire T93;
  wire[1:0] T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[1:0] T98;
  wire[1:0] T99;
  wire[7:0] T100;
  wire[3:0] T101;
  wire[1:0] T102;
  wire T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[3:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire[3:0] T110;
  wire[1:0] T111;
  wire[7:0] T112;
  wire[3:0] T113;
  wire[1:0] T114;
  wire T115;
  wire[1:0] T116;
  wire T117;
  wire[3:0] T118;
  wire[1:0] T119;
  wire[7:0] T120;
  wire[3:0] T121;
  wire[1:0] T122;
  wire T123;
  wire[1:0] T124;
  wire T125;
  wire[3:0] T126;
  wire[1:0] T127;
  wire[3:0] T128;
  wire[2:0] T129;
  wire[7:0] T130;
  wire[3:0] T131;
  wire[1:0] T132;
  wire T133;
  wire[1:0] T134;
  wire T135;
  wire T136;
  wire[3:0] T137;
  wire[2:0] T138;
  wire[7:0] T139;
  wire[3:0] T140;
  wire[1:0] T141;
  wire T142;
  wire[1:0] T143;
  wire T144;
  wire T145;
  wire[3:0] T146;
  wire[2:0] T147;
  wire[3:0] T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire[7:0] T151;
  wire[3:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[1:0] T160;
  wire[1:0] T161;
  wire[7:0] T162;
  wire[3:0] T163;
  wire[1:0] T164;
  wire T165;
  wire T166;
  wire[1:0] T167;
  wire T168;
  wire T169;
  wire[3:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire[3:0] T173;
  wire[1:0] T174;
  wire[1:0] T175;
  wire[7:0] T176;
  wire[3:0] T177;
  wire[1:0] T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire[3:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire[7:0] T187;
  wire[3:0] T188;
  wire[1:0] T189;
  wire T190;
  wire T191;
  wire[1:0] T192;
  wire T193;
  wire T194;
  wire[3:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[3:0] T198;
  wire[1:0] T199;
  wire[1:0] T200;
  wire[7:0] T201;
  wire[3:0] T202;
  wire[1:0] T203;
  wire T204;
  wire T205;
  wire[1:0] T206;
  wire T207;
  wire T208;
  wire[3:0] T209;
  wire[1:0] T210;
  wire[1:0] T211;
  wire[7:0] T212;
  wire[3:0] T213;
  wire[1:0] T214;
  wire T215;
  wire T216;
  wire[1:0] T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[1:0] T221;
  wire[1:0] T222;
  wire[3:0] T223;
  wire[1:0] T224;
  wire[1:0] T225;
  wire[7:0] T226;
  wire[3:0] T227;
  wire[1:0] T228;
  wire T229;
  wire T230;
  wire[1:0] T231;
  wire T232;
  wire T233;
  wire[3:0] T234;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[7:0] T237;
  wire[3:0] T238;
  wire[1:0] T239;
  wire T240;
  wire T241;
  wire[1:0] T242;
  wire T243;
  wire T244;
  wire[3:0] T245;
  wire[1:0] T246;
  wire[1:0] T247;
  wire[3:0] T248;
  wire[1:0] T249;
  wire[7:0] T250;
  wire[3:0] T251;
  wire[1:0] T252;
  wire T253;
  wire T254;
  wire[1:0] T255;
  wire T256;
  wire[3:0] T257;
  wire[1:0] T258;
  wire[7:0] T259;
  wire[3:0] T260;
  wire[1:0] T261;
  wire T262;
  wire T263;
  wire[1:0] T264;
  wire T265;
  wire[3:0] T266;
  wire[1:0] T267;
  wire[3:0] T268;
  wire[2:0] T269;
  wire[7:0] T270;
  wire[3:0] T271;
  wire[1:0] T272;
  wire T273;
  wire[1:0] T274;
  wire T275;
  wire T276;
  wire[3:0] T277;
  wire[2:0] T278;
  wire[7:0] T279;
  wire[3:0] T280;
  wire[1:0] T281;
  wire T282;
  wire[1:0] T283;
  wire T284;
  wire T285;
  wire[3:0] T286;
  wire[2:0] T287;
  wire[3:0] T288;
  wire[1:0] T289;
  wire[1:0] T290;
  wire[7:0] T291;
  wire[3:0] T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire[1:0] T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[7:0] T302;
  wire[3:0] T303;
  wire[1:0] T304;
  wire T305;
  wire T306;
  wire[1:0] T307;
  wire T308;
  wire T309;
  wire[3:0] T310;
  wire[1:0] T311;
  wire[1:0] T312;
  wire[3:0] T313;
  wire[1:0] T314;
  wire[1:0] T315;
  wire[7:0] T316;
  wire[3:0] T317;
  wire[1:0] T318;
  wire T319;
  wire T320;
  wire[1:0] T321;
  wire T322;
  wire T323;
  wire[3:0] T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[7:0] T327;
  wire[3:0] T328;
  wire[1:0] T329;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire T333;
  wire T334;
  wire[3:0] T335;
  wire[1:0] T336;
  wire[1:0] T337;
  wire[3:0] T338;
  wire[1:0] T339;
  wire[1:0] T340;
  wire[7:0] T341;
  wire[3:0] T342;
  wire[1:0] T343;
  wire T344;
  wire T345;
  wire[1:0] T346;
  wire T347;
  wire T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire[1:0] T351;
  wire[7:0] T352;
  wire[3:0] T353;
  wire[1:0] T354;
  wire T355;
  wire T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire[3:0] T360;
  wire[1:0] T361;
  wire[1:0] T362;
  wire[3:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[7:0] T366;
  wire[3:0] T367;
  wire[1:0] T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire T372;
  wire T373;
  wire[3:0] T374;
  wire[1:0] T375;
  wire[1:0] T376;
  wire[7:0] T377;
  wire[3:0] T378;
  wire[1:0] T379;
  wire T380;
  wire T381;
  wire[1:0] T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[3:0] T388;
  wire[1:0] T389;
  wire[7:0] T390;
  wire[3:0] T391;
  wire[1:0] T392;
  wire T393;
  wire T394;
  wire[1:0] T395;
  wire T396;
  wire[3:0] T397;
  wire[1:0] T398;
  wire[7:0] T399;
  wire[3:0] T400;
  wire[1:0] T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire T405;
  wire[3:0] T406;
  wire[1:0] T407;
  wire[3:0] T408;
  wire[2:0] T409;
  wire[7:0] T410;
  wire[3:0] T411;
  wire[1:0] T412;
  wire T413;
  wire[1:0] T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[2:0] T418;
  wire[7:0] T419;
  wire[3:0] T420;
  wire[1:0] T421;
  wire T422;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire[3:0] T426;
  wire[2:0] T427;
  wire[3:0] T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire[7:0] T431;
  wire[3:0] T432;
  wire[1:0] T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire T437;
  wire T438;
  wire[3:0] T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire[7:0] T442;
  wire[3:0] T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire[1:0] T447;
  wire T448;
  wire T449;
  wire[3:0] T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[3:0] T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire[7:0] T456;
  wire[3:0] T457;
  wire[1:0] T458;
  wire T459;
  wire T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire[3:0] T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[7:0] T467;
  wire[3:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire T473;
  wire T474;
  wire[3:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[3:0] T478;
  wire[1:0] T479;
  wire[1:0] T480;
  wire[7:0] T481;
  wire[3:0] T482;
  wire[1:0] T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[1:0] T490;
  wire[1:0] T491;
  wire[7:0] T492;
  wire[3:0] T493;
  wire[1:0] T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire T498;
  wire T499;
  wire[3:0] T500;
  wire[1:0] T501;
  wire[1:0] T502;
  wire[3:0] T503;
  wire[1:0] T504;
  wire[1:0] T505;
  wire[7:0] T506;
  wire[3:0] T507;
  wire[1:0] T508;
  wire T509;
  wire T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire[3:0] T514;
  wire[1:0] T515;
  wire[1:0] T516;
  wire[7:0] T517;
  wire[3:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire[1:0] T522;
  wire T523;
  wire T524;
  wire[3:0] T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire[3:0] T528;
  wire[1:0] T529;
  wire[7:0] T530;
  wire[3:0] T531;
  wire[1:0] T532;
  wire T533;
  wire T534;
  wire[1:0] T535;
  wire T536;
  wire[3:0] T537;
  wire[1:0] T538;
  wire[7:0] T539;
  wire[3:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire T545;
  wire[3:0] T546;
  wire[1:0] T547;
  wire[3:0] T548;
  wire[2:0] T549;
  wire[7:0] T550;
  wire[3:0] T551;
  wire[1:0] T552;
  wire T553;
  wire[1:0] T554;
  wire T555;
  wire T556;
  wire[3:0] T557;
  wire[2:0] T558;
  wire[7:0] T559;
  wire[3:0] T560;
  wire[1:0] T561;
  wire T562;
  wire[1:0] T563;
  wire T564;
  wire T565;
  wire[3:0] T566;
  wire[2:0] T567;
  wire[3:0] T568;
  wire[1:0] T569;
  wire[1:0] T570;
  wire[7:0] T571;
  wire[3:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire[1:0] T576;
  wire T577;
  wire T578;
  wire[3:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[7:0] T582;
  wire[3:0] T583;
  wire[1:0] T584;
  wire T585;
  wire T586;
  wire[1:0] T587;
  wire T588;
  wire T589;
  wire[3:0] T590;
  wire[1:0] T591;
  wire[1:0] T592;
  wire[3:0] T593;
  wire[1:0] T594;
  wire[1:0] T595;
  wire[7:0] T596;
  wire[3:0] T597;
  wire[1:0] T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire T602;
  wire T603;
  wire[3:0] T604;
  wire[1:0] T605;
  wire[1:0] T606;
  wire[7:0] T607;
  wire[3:0] T608;
  wire[1:0] T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire T613;
  wire T614;
  wire[3:0] T615;
  wire[1:0] T616;
  wire[1:0] T617;
  wire[3:0] T618;
  wire[1:0] T619;
  wire[1:0] T620;
  wire[7:0] T621;
  wire[3:0] T622;
  wire[1:0] T623;
  wire T624;
  wire T625;
  wire[1:0] T626;
  wire T627;
  wire T628;
  wire[3:0] T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire[7:0] T632;
  wire[3:0] T633;
  wire[1:0] T634;
  wire T635;
  wire T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire[3:0] T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[3:0] T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire[7:0] T646;
  wire[3:0] T647;
  wire[1:0] T648;
  wire T649;
  wire T650;
  wire[1:0] T651;
  wire T652;
  wire T653;
  wire[3:0] T654;
  wire[1:0] T655;
  wire[1:0] T656;
  wire[7:0] T657;
  wire[3:0] T658;
  wire[1:0] T659;
  wire T660;
  wire T661;
  wire[1:0] T662;
  wire T663;
  wire T664;
  wire[3:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[3:0] T668;
  wire[1:0] T669;
  wire[7:0] T670;
  wire[3:0] T671;
  wire[1:0] T672;
  wire T673;
  wire T674;
  wire[1:0] T675;
  wire T676;
  wire[3:0] T677;
  wire[1:0] T678;
  wire[7:0] T679;
  wire[3:0] T680;
  wire[1:0] T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire T685;
  wire[3:0] T686;
  wire[1:0] T687;
  wire[3:0] T688;
  wire[7:0] T689;
  wire[2:0] T690;
  wire[1:0] T691;
  wire T692;
  wire[4:0] T693;
  wire[3:0] T694;
  wire T695;
  wire[7:0] T696;
  wire[2:0] T697;
  wire[1:0] T698;
  wire T699;
  wire[4:0] T700;
  wire[3:0] T701;
  wire T702;
  wire[3:0] T703;
  wire[2:0] T704;
  wire[7:0] T705;
  wire[3:0] T706;
  wire[1:0] T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire T711;
  wire[3:0] T712;
  wire[2:0] T713;
  wire[7:0] T714;
  wire[3:0] T715;
  wire[1:0] T716;
  wire T717;
  wire T718;
  wire[1:0] T719;
  wire T720;
  wire[3:0] T721;
  wire[2:0] T722;
  wire[3:0] T723;
  wire[2:0] T724;
  wire[7:0] T725;
  wire[3:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire[1:0] T730;
  wire T731;
  wire[3:0] T732;
  wire[2:0] T733;
  wire[7:0] T734;
  wire[3:0] T735;
  wire[1:0] T736;
  wire T737;
  wire T738;
  wire[1:0] T739;
  wire T740;
  wire[3:0] T741;
  wire[2:0] T742;
  wire[3:0] T743;
  wire[2:0] T744;
  wire[7:0] T745;
  wire[3:0] T746;
  wire[1:0] T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire T751;
  wire[3:0] T752;
  wire[2:0] T753;
  wire[7:0] T754;
  wire[3:0] T755;
  wire[1:0] T756;
  wire T757;
  wire T758;
  wire[1:0] T759;
  wire T760;
  wire[3:0] T761;
  wire[2:0] T762;
  wire[3:0] T763;
  wire[2:0] T764;
  wire[7:0] T765;
  wire[3:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire[1:0] T770;
  wire T771;
  wire[3:0] T772;
  wire[2:0] T773;
  wire[7:0] T774;
  wire[3:0] T775;
  wire[1:0] T776;
  wire T777;
  wire T778;
  wire[1:0] T779;
  wire T780;
  wire[3:0] T781;
  wire[2:0] T782;
  wire[3:0] T783;
  wire[7:0] T784;
  wire[2:0] T785;
  wire[1:0] T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire[1:0] T790;
  wire[7:0] T791;
  wire[2:0] T792;
  wire[1:0] T793;
  wire T794;
  wire T795;
  wire[4:0] T796;
  wire[1:0] T797;
  wire[3:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire[1:0] T802;
  wire T803;
  wire T804;
  wire[3:0] T805;
  wire[1:0] T806;
  wire T807;
  wire T808;
  wire[1:0] T809;
  wire T810;
  wire T811;
  wire[3:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire[1:0] T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[1:0] T820;
  wire T821;
  wire T822;
  wire[1:0] T823;
  wire T824;
  wire T825;
  wire[3:0] T826;
  wire[1:0] T827;
  wire T828;
  wire T829;
  wire[1:0] T830;
  wire T831;
  wire T832;
  wire[3:0] T833;
  wire[1:0] T834;
  wire T835;
  wire T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire[3:0] T840;
  wire[1:0] T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire T845;
  wire T846;
  wire[3:0] T847;
  wire[1:0] T848;
  wire T849;
  wire T850;
  wire[1:0] T851;
  wire T852;
  wire T853;
  wire[3:0] T854;
  wire[1:0] T855;
  wire T856;
  wire T857;
  wire[1:0] T858;
  wire T859;
  wire T860;
  wire[3:0] T861;
  wire[1:0] T862;
  wire T863;
  wire T864;
  wire[1:0] T865;
  wire T866;
  wire T867;
  wire[3:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire[1:0] T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[1:0] T876;
  wire T877;
  wire T878;
  wire[1:0] T879;
  wire T880;
  wire T881;
  wire[3:0] T882;
  wire[1:0] T883;
  wire T884;
  wire T885;
  wire[1:0] T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[1:0] T890;
  wire T891;
  wire T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire[3:0] T896;
  wire[1:0] T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire T901;
  wire T902;
  wire[3:0] T903;
  wire[1:0] T904;
  wire T905;
  wire T906;
  wire[1:0] T907;
  wire T908;
  wire T909;
  wire[3:0] T910;
  wire[1:0] T911;
  wire T912;
  wire T913;
  wire[1:0] T914;
  wire T915;
  wire T916;
  wire[3:0] T917;
  wire[1:0] T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire T922;
  wire T923;
  wire[3:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire[1:0] T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[1:0] T932;
  wire T933;
  wire T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire[3:0] T938;
  wire[1:0] T939;
  wire T940;
  wire T941;
  wire[1:0] T942;
  wire T943;
  wire T944;
  wire[3:0] T945;
  wire[1:0] T946;
  wire T947;
  wire T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire[3:0] T952;
  wire[1:0] T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire T957;
  wire T958;
  wire[3:0] T959;
  wire[1:0] T960;
  wire T961;
  wire T962;
  wire[1:0] T963;
  wire T964;
  wire T965;
  wire[3:0] T966;
  wire[1:0] T967;
  wire T968;
  wire T969;
  wire[1:0] T970;
  wire T971;
  wire T972;
  wire[3:0] T973;
  wire[1:0] T974;
  wire T975;
  wire T976;
  wire[1:0] T977;
  wire T978;
  wire T979;
  wire[3:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire[1:0] T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[1:0] T988;
  wire T989;
  wire T990;
  wire[1:0] T991;
  wire T992;
  wire T993;
  wire[3:0] T994;
  wire[1:0] T995;
  wire T996;
  wire T997;
  wire[1:0] T998;
  wire T999;
  wire T1000;
  wire[3:0] T1001;
  wire[1:0] T1002;
  wire T1003;
  wire T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire[3:0] T1008;
  wire[1:0] T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire T1013;
  wire T1014;
  wire[3:0] T1015;
  wire[1:0] T1016;
  wire T1017;
  wire T1018;
  wire[1:0] T1019;
  wire T1020;
  wire T1021;
  wire[3:0] T1022;
  wire[1:0] T1023;
  wire T1024;
  wire T1025;
  wire[1:0] T1026;
  wire T1027;
  wire T1028;
  wire[3:0] T1029;
  wire[1:0] T1030;
  wire T1031;
  wire T1032;
  wire[1:0] T1033;
  wire T1034;
  wire T1035;
  wire[3:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire[1:0] T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[1:0] T1044;
  wire T1045;
  wire T1046;
  wire[1:0] T1047;
  wire T1048;
  wire T1049;
  wire[3:0] T1050;
  wire[1:0] T1051;
  wire T1052;
  wire T1053;
  wire[1:0] T1054;
  wire T1055;
  wire T1056;
  wire[3:0] T1057;
  wire[1:0] T1058;
  wire T1059;
  wire T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire[3:0] T1064;
  wire[1:0] T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire T1069;
  wire T1070;
  wire[3:0] T1071;
  wire[1:0] T1072;
  wire T1073;
  wire T1074;
  wire[1:0] T1075;
  wire T1076;
  wire T1077;
  wire[3:0] T1078;
  wire[1:0] T1079;
  wire T1080;
  wire T1081;
  wire[1:0] T1082;
  wire T1083;
  wire T1084;
  wire[3:0] T1085;
  wire[1:0] T1086;
  wire T1087;
  wire T1088;
  wire[1:0] T1089;
  wire T1090;
  wire T1091;
  wire[3:0] T1092;
  wire[1:0] T1093;
  wire T1094;
  wire T1095;
  wire[1:0] T1096;
  wire T1097;
  wire T1098;
  wire[3:0] T1099;
  wire[1:0] T1100;
  wire T1101;
  wire T1102;
  wire[1:0] T1103;
  wire T1104;
  wire T1105;
  wire[3:0] T1106;
  wire[1:0] T1107;
  wire T1108;
  wire T1109;
  wire[1:0] T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[1:0] T1114;
  wire T1115;
  wire T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire[3:0] T1120;
  wire[1:0] T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[1:0] T1128;
  wire T1129;
  wire T1130;
  wire[1:0] T1131;
  wire T1132;
  wire T1133;
  wire[3:0] T1134;
  wire[1:0] T1135;
  wire T1136;
  wire T1137;
  wire[1:0] T1138;
  wire T1139;
  wire T1140;
  wire[3:0] T1141;
  wire[1:0] T1142;
  wire T1143;
  wire T1144;
  wire[1:0] T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire[32:0] CU_io_out;
  wire CU_io_enqRdy;
  wire CU_io_deqValid;
  wire CU_io_enqRdyOut;
  wire[32:0] CU_1_io_out;
  wire CU_1_io_enqRdy;
  wire CU_1_io_deqValid;
  wire CU_1_io_enqRdyOut;
  wire[32:0] CU_2_io_out;
  wire CU_2_io_enqRdy;
  wire CU_2_io_deqValid;
  wire CU_2_io_enqRdyOut;
  wire[32:0] CU_3_io_out;
  wire CU_3_io_enqRdy;
  wire CU_3_io_deqValid;
  wire CU_3_io_enqRdyOut;
  wire[32:0] CU_4_io_out;
  wire CU_4_io_enqRdy;
  wire CU_4_io_deqValid;
  wire CU_4_io_enqRdyOut;
  wire[32:0] CU_5_io_out;
  wire CU_5_io_enqRdy;
  wire CU_5_io_deqValid;
  wire CU_5_io_enqRdyOut;
  wire[32:0] CU_6_io_out;
  wire CU_6_io_enqRdy;
  wire CU_6_io_deqValid;
  wire CU_6_io_enqRdyOut;
  wire[32:0] CU_7_io_out;
  wire CU_7_io_enqRdy;
  wire CU_7_io_deqValid;
  wire CU_7_io_enqRdyOut;
  wire[32:0] CU_8_io_out;
  wire CU_8_io_enqRdy;
  wire CU_8_io_deqValid;
  wire CU_8_io_enqRdyOut;
  wire[32:0] CU_9_io_out;
  wire CU_9_io_enqRdy;
  wire CU_9_io_deqValid;
  wire CU_9_io_enqRdyOut;
  wire[32:0] CU_10_io_out;
  wire CU_10_io_enqRdy;
  wire CU_10_io_deqValid;
  wire CU_10_io_enqRdyOut;
  wire[32:0] CU_11_io_out;
  wire CU_11_io_enqRdy;
  wire CU_11_io_deqValid;
  wire CU_11_io_enqRdyOut;
  wire[32:0] CU_12_io_out;
  wire CU_12_io_enqRdy;
  wire CU_12_io_deqValid;
  wire CU_12_io_enqRdyOut;
  wire[32:0] CU_13_io_out;
  wire CU_13_io_enqRdy;
  wire CU_13_io_deqValid;
  wire CU_13_io_enqRdyOut;
  wire[32:0] CU_14_io_out;
  wire CU_14_io_enqRdy;
  wire CU_14_io_deqValid;
  wire CU_14_io_enqRdyOut;
  wire[32:0] CU_15_io_out;
  wire CU_15_io_enqRdy;
  wire CU_15_io_deqValid;
  wire CU_15_io_enqRdyOut;
  wire[32:0] CU_16_io_out;
  wire CU_16_io_enqRdy;
  wire CU_16_io_deqValid;
  wire CU_16_io_enqRdyOut;
  wire[32:0] CU_17_io_out;
  wire CU_17_io_enqRdy;
  wire CU_17_io_deqValid;
  wire CU_17_io_enqRdyOut;
  wire[32:0] CU_18_io_out;
  wire CU_18_io_enqRdy;
  wire CU_18_io_deqValid;
  wire CU_18_io_enqRdyOut;
  wire[32:0] CU_19_io_out;
  wire CU_19_io_enqRdy;
  wire CU_19_io_deqValid;
  wire CU_19_io_enqRdyOut;
  wire[32:0] CU_20_io_out;
  wire CU_20_io_enqRdy;
  wire CU_20_io_deqValid;
  wire CU_20_io_enqRdyOut;
  wire[32:0] CU_21_io_out;
  wire CU_21_io_enqRdy;
  wire CU_21_io_deqValid;
  wire CU_21_io_enqRdyOut;
  wire[32:0] CU_22_io_out;
  wire CU_22_io_enqRdy;
  wire CU_22_io_deqValid;
  wire CU_22_io_enqRdyOut;
  wire[32:0] CU_23_io_out;
  wire CU_23_io_enqRdy;
  wire CU_23_io_deqValid;
  wire CU_23_io_enqRdyOut;
  wire[32:0] CU_24_io_out;
  wire CU_24_io_enqRdy;
  wire CU_24_io_deqValid;
  wire CU_24_io_enqRdyOut;
  wire[32:0] Switch_io_outPort_4;
  wire[32:0] Switch_io_outPort_3;
  wire[32:0] Switch_io_outPort_1;
  wire[32:0] Switch_io_outPort_0;
  wire[7:0] Switch_io_deqValid;
  wire[7:0] Switch_io_enqRdy;
  wire[23:0] Switch_io_outCUConfig;
  wire[32:0] Switch_1_io_outPort_7;
  wire[32:0] Switch_1_io_outPort_4;
  wire[32:0] Switch_1_io_outPort_3;
  wire[32:0] Switch_1_io_outPort_2;
  wire[32:0] Switch_1_io_outPort_1;
  wire[32:0] Switch_1_io_outPort_0;
  wire[7:0] Switch_1_io_deqValid;
  wire[7:0] Switch_1_io_enqRdy;
  wire[23:0] Switch_1_io_outCUConfig;
  wire Switch_1_io_enqOR;
  wire[32:0] Switch_2_io_outPort_7;
  wire[32:0] Switch_2_io_outPort_4;
  wire[32:0] Switch_2_io_outPort_3;
  wire[32:0] Switch_2_io_outPort_2;
  wire[32:0] Switch_2_io_outPort_1;
  wire[32:0] Switch_2_io_outPort_0;
  wire[7:0] Switch_2_io_deqValid;
  wire[7:0] Switch_2_io_enqRdy;
  wire[23:0] Switch_2_io_outCUConfig;
  wire Switch_2_io_enqOR;
  wire[32:0] Switch_3_io_outPort_7;
  wire[32:0] Switch_3_io_outPort_4;
  wire[32:0] Switch_3_io_outPort_3;
  wire[32:0] Switch_3_io_outPort_2;
  wire[32:0] Switch_3_io_outPort_1;
  wire[32:0] Switch_3_io_outPort_0;
  wire[7:0] Switch_3_io_deqValid;
  wire[7:0] Switch_3_io_enqRdy;
  wire[23:0] Switch_3_io_outCUConfig;
  wire Switch_3_io_enqOR;
  wire[32:0] Switch_4_io_outPort_7;
  wire[32:0] Switch_4_io_outPort_4;
  wire[32:0] Switch_4_io_outPort_3;
  wire[32:0] Switch_4_io_outPort_2;
  wire[32:0] Switch_4_io_outPort_1;
  wire[32:0] Switch_4_io_outPort_0;
  wire[7:0] Switch_4_io_deqValid;
  wire[7:0] Switch_4_io_enqRdy;
  wire[23:0] Switch_4_io_outCUConfig;
  wire Switch_4_io_enqOR;
  wire[32:0] Switch_5_io_outPort_7;
  wire[32:0] Switch_5_io_outPort_3;
  wire[32:0] Switch_5_io_outPort_1;
  wire[32:0] Switch_5_io_outPort_0;
  wire[7:0] Switch_5_io_deqValid;
  wire[7:0] Switch_5_io_enqRdy;
  wire Switch_5_io_enqOR;
  wire[32:0] Switch_6_io_outPort_5;
  wire[32:0] Switch_6_io_outPort_4;
  wire[32:0] Switch_6_io_outPort_3;
  wire[32:0] Switch_6_io_outPort_2;
  wire[32:0] Switch_6_io_outPort_1;
  wire[32:0] Switch_6_io_outPort_0;
  wire[7:0] Switch_6_io_deqValid;
  wire[7:0] Switch_6_io_enqRdy;
  wire[23:0] Switch_6_io_outCUConfig;
  wire[32:0] Switch_7_io_outPort_7;
  wire[32:0] Switch_7_io_outPort_6;
  wire[32:0] Switch_7_io_outPort_5;
  wire[32:0] Switch_7_io_outPort_4;
  wire[32:0] Switch_7_io_outPort_3;
  wire[32:0] Switch_7_io_outPort_2;
  wire[32:0] Switch_7_io_outPort_1;
  wire[32:0] Switch_7_io_outPort_0;
  wire[7:0] Switch_7_io_deqValid;
  wire[7:0] Switch_7_io_enqRdy;
  wire[23:0] Switch_7_io_outCUConfig;
  wire Switch_7_io_enqOR;
  wire[32:0] Switch_8_io_outPort_7;
  wire[32:0] Switch_8_io_outPort_6;
  wire[32:0] Switch_8_io_outPort_5;
  wire[32:0] Switch_8_io_outPort_4;
  wire[32:0] Switch_8_io_outPort_3;
  wire[32:0] Switch_8_io_outPort_2;
  wire[32:0] Switch_8_io_outPort_1;
  wire[32:0] Switch_8_io_outPort_0;
  wire[7:0] Switch_8_io_deqValid;
  wire[7:0] Switch_8_io_enqRdy;
  wire[23:0] Switch_8_io_outCUConfig;
  wire Switch_8_io_enqOR;
  wire[32:0] Switch_9_io_outPort_7;
  wire[32:0] Switch_9_io_outPort_6;
  wire[32:0] Switch_9_io_outPort_5;
  wire[32:0] Switch_9_io_outPort_4;
  wire[32:0] Switch_9_io_outPort_3;
  wire[32:0] Switch_9_io_outPort_2;
  wire[32:0] Switch_9_io_outPort_1;
  wire[32:0] Switch_9_io_outPort_0;
  wire[7:0] Switch_9_io_deqValid;
  wire[7:0] Switch_9_io_enqRdy;
  wire[23:0] Switch_9_io_outCUConfig;
  wire Switch_9_io_enqOR;
  wire[32:0] Switch_10_io_outPort_7;
  wire[32:0] Switch_10_io_outPort_6;
  wire[32:0] Switch_10_io_outPort_5;
  wire[32:0] Switch_10_io_outPort_4;
  wire[32:0] Switch_10_io_outPort_3;
  wire[32:0] Switch_10_io_outPort_2;
  wire[32:0] Switch_10_io_outPort_1;
  wire[32:0] Switch_10_io_outPort_0;
  wire[7:0] Switch_10_io_deqValid;
  wire[7:0] Switch_10_io_enqRdy;
  wire[23:0] Switch_10_io_outCUConfig;
  wire Switch_10_io_enqOR;
  wire[32:0] Switch_11_io_outPort_7;
  wire[32:0] Switch_11_io_outPort_6;
  wire[32:0] Switch_11_io_outPort_3;
  wire[32:0] Switch_11_io_outPort_2;
  wire[32:0] Switch_11_io_outPort_1;
  wire[32:0] Switch_11_io_outPort_0;
  wire[7:0] Switch_11_io_deqValid;
  wire[7:0] Switch_11_io_enqRdy;
  wire Switch_11_io_enqOR;
  wire[32:0] Switch_12_io_outPort_5;
  wire[32:0] Switch_12_io_outPort_4;
  wire[32:0] Switch_12_io_outPort_3;
  wire[32:0] Switch_12_io_outPort_2;
  wire[32:0] Switch_12_io_outPort_1;
  wire[32:0] Switch_12_io_outPort_0;
  wire[7:0] Switch_12_io_deqValid;
  wire[7:0] Switch_12_io_enqRdy;
  wire[23:0] Switch_12_io_outCUConfig;
  wire[32:0] Switch_13_io_outPort_7;
  wire[32:0] Switch_13_io_outPort_6;
  wire[32:0] Switch_13_io_outPort_5;
  wire[32:0] Switch_13_io_outPort_4;
  wire[32:0] Switch_13_io_outPort_3;
  wire[32:0] Switch_13_io_outPort_2;
  wire[32:0] Switch_13_io_outPort_1;
  wire[32:0] Switch_13_io_outPort_0;
  wire[7:0] Switch_13_io_deqValid;
  wire[7:0] Switch_13_io_enqRdy;
  wire[23:0] Switch_13_io_outCUConfig;
  wire Switch_13_io_enqOR;
  wire[32:0] Switch_14_io_outPort_7;
  wire[32:0] Switch_14_io_outPort_6;
  wire[32:0] Switch_14_io_outPort_5;
  wire[32:0] Switch_14_io_outPort_4;
  wire[32:0] Switch_14_io_outPort_3;
  wire[32:0] Switch_14_io_outPort_2;
  wire[32:0] Switch_14_io_outPort_1;
  wire[32:0] Switch_14_io_outPort_0;
  wire[7:0] Switch_14_io_deqValid;
  wire[7:0] Switch_14_io_enqRdy;
  wire[23:0] Switch_14_io_outCUConfig;
  wire Switch_14_io_enqOR;
  wire[32:0] Switch_15_io_outPort_7;
  wire[32:0] Switch_15_io_outPort_6;
  wire[32:0] Switch_15_io_outPort_5;
  wire[32:0] Switch_15_io_outPort_4;
  wire[32:0] Switch_15_io_outPort_3;
  wire[32:0] Switch_15_io_outPort_2;
  wire[32:0] Switch_15_io_outPort_1;
  wire[32:0] Switch_15_io_outPort_0;
  wire[7:0] Switch_15_io_deqValid;
  wire[7:0] Switch_15_io_enqRdy;
  wire[23:0] Switch_15_io_outCUConfig;
  wire Switch_15_io_enqOR;
  wire[32:0] Switch_16_io_outPort_7;
  wire[32:0] Switch_16_io_outPort_6;
  wire[32:0] Switch_16_io_outPort_5;
  wire[32:0] Switch_16_io_outPort_4;
  wire[32:0] Switch_16_io_outPort_3;
  wire[32:0] Switch_16_io_outPort_2;
  wire[32:0] Switch_16_io_outPort_1;
  wire[32:0] Switch_16_io_outPort_0;
  wire[7:0] Switch_16_io_deqValid;
  wire[7:0] Switch_16_io_enqRdy;
  wire[23:0] Switch_16_io_outCUConfig;
  wire Switch_16_io_enqOR;
  wire[32:0] Switch_17_io_outPort_7;
  wire[32:0] Switch_17_io_outPort_6;
  wire[32:0] Switch_17_io_outPort_3;
  wire[32:0] Switch_17_io_outPort_2;
  wire[32:0] Switch_17_io_outPort_1;
  wire[32:0] Switch_17_io_outPort_0;
  wire[7:0] Switch_17_io_deqValid;
  wire[7:0] Switch_17_io_enqRdy;
  wire Switch_17_io_enqOR;
  wire[32:0] Switch_18_io_outPort_5;
  wire[32:0] Switch_18_io_outPort_4;
  wire[32:0] Switch_18_io_outPort_3;
  wire[32:0] Switch_18_io_outPort_2;
  wire[32:0] Switch_18_io_outPort_1;
  wire[32:0] Switch_18_io_outPort_0;
  wire[7:0] Switch_18_io_deqValid;
  wire[7:0] Switch_18_io_enqRdy;
  wire[23:0] Switch_18_io_outCUConfig;
  wire[32:0] Switch_19_io_outPort_7;
  wire[32:0] Switch_19_io_outPort_6;
  wire[32:0] Switch_19_io_outPort_5;
  wire[32:0] Switch_19_io_outPort_4;
  wire[32:0] Switch_19_io_outPort_3;
  wire[32:0] Switch_19_io_outPort_2;
  wire[32:0] Switch_19_io_outPort_1;
  wire[32:0] Switch_19_io_outPort_0;
  wire[7:0] Switch_19_io_deqValid;
  wire[7:0] Switch_19_io_enqRdy;
  wire[23:0] Switch_19_io_outCUConfig;
  wire Switch_19_io_enqOR;
  wire[32:0] Switch_20_io_outPort_7;
  wire[32:0] Switch_20_io_outPort_6;
  wire[32:0] Switch_20_io_outPort_5;
  wire[32:0] Switch_20_io_outPort_4;
  wire[32:0] Switch_20_io_outPort_3;
  wire[32:0] Switch_20_io_outPort_2;
  wire[32:0] Switch_20_io_outPort_1;
  wire[32:0] Switch_20_io_outPort_0;
  wire[7:0] Switch_20_io_deqValid;
  wire[7:0] Switch_20_io_enqRdy;
  wire[23:0] Switch_20_io_outCUConfig;
  wire Switch_20_io_enqOR;
  wire[32:0] Switch_21_io_outPort_7;
  wire[32:0] Switch_21_io_outPort_6;
  wire[32:0] Switch_21_io_outPort_5;
  wire[32:0] Switch_21_io_outPort_4;
  wire[32:0] Switch_21_io_outPort_3;
  wire[32:0] Switch_21_io_outPort_2;
  wire[32:0] Switch_21_io_outPort_1;
  wire[32:0] Switch_21_io_outPort_0;
  wire[7:0] Switch_21_io_deqValid;
  wire[7:0] Switch_21_io_enqRdy;
  wire[23:0] Switch_21_io_outCUConfig;
  wire Switch_21_io_enqOR;
  wire[32:0] Switch_22_io_outPort_7;
  wire[32:0] Switch_22_io_outPort_6;
  wire[32:0] Switch_22_io_outPort_5;
  wire[32:0] Switch_22_io_outPort_4;
  wire[32:0] Switch_22_io_outPort_3;
  wire[32:0] Switch_22_io_outPort_2;
  wire[32:0] Switch_22_io_outPort_1;
  wire[32:0] Switch_22_io_outPort_0;
  wire[7:0] Switch_22_io_deqValid;
  wire[7:0] Switch_22_io_enqRdy;
  wire[23:0] Switch_22_io_outCUConfig;
  wire Switch_22_io_enqOR;
  wire[32:0] Switch_23_io_outPort_7;
  wire[32:0] Switch_23_io_outPort_6;
  wire[32:0] Switch_23_io_outPort_3;
  wire[32:0] Switch_23_io_outPort_2;
  wire[32:0] Switch_23_io_outPort_1;
  wire[32:0] Switch_23_io_outPort_0;
  wire[7:0] Switch_23_io_deqValid;
  wire[7:0] Switch_23_io_enqRdy;
  wire Switch_23_io_enqOR;
  wire[32:0] Switch_24_io_outPort_5;
  wire[32:0] Switch_24_io_outPort_4;
  wire[32:0] Switch_24_io_outPort_3;
  wire[32:0] Switch_24_io_outPort_2;
  wire[32:0] Switch_24_io_outPort_1;
  wire[32:0] Switch_24_io_outPort_0;
  wire[7:0] Switch_24_io_deqValid;
  wire[7:0] Switch_24_io_enqRdy;
  wire[23:0] Switch_24_io_outCUConfig;
  wire[32:0] Switch_25_io_outPort_7;
  wire[32:0] Switch_25_io_outPort_6;
  wire[32:0] Switch_25_io_outPort_5;
  wire[32:0] Switch_25_io_outPort_4;
  wire[32:0] Switch_25_io_outPort_3;
  wire[32:0] Switch_25_io_outPort_2;
  wire[32:0] Switch_25_io_outPort_1;
  wire[32:0] Switch_25_io_outPort_0;
  wire[7:0] Switch_25_io_deqValid;
  wire[7:0] Switch_25_io_enqRdy;
  wire[23:0] Switch_25_io_outCUConfig;
  wire Switch_25_io_enqOR;
  wire[32:0] Switch_26_io_outPort_7;
  wire[32:0] Switch_26_io_outPort_6;
  wire[32:0] Switch_26_io_outPort_5;
  wire[32:0] Switch_26_io_outPort_4;
  wire[32:0] Switch_26_io_outPort_3;
  wire[32:0] Switch_26_io_outPort_2;
  wire[32:0] Switch_26_io_outPort_1;
  wire[32:0] Switch_26_io_outPort_0;
  wire[7:0] Switch_26_io_deqValid;
  wire[7:0] Switch_26_io_enqRdy;
  wire[23:0] Switch_26_io_outCUConfig;
  wire Switch_26_io_enqOR;
  wire[32:0] Switch_27_io_outPort_7;
  wire[32:0] Switch_27_io_outPort_6;
  wire[32:0] Switch_27_io_outPort_5;
  wire[32:0] Switch_27_io_outPort_4;
  wire[32:0] Switch_27_io_outPort_3;
  wire[32:0] Switch_27_io_outPort_2;
  wire[32:0] Switch_27_io_outPort_1;
  wire[32:0] Switch_27_io_outPort_0;
  wire[7:0] Switch_27_io_deqValid;
  wire[7:0] Switch_27_io_enqRdy;
  wire[23:0] Switch_27_io_outCUConfig;
  wire Switch_27_io_enqOR;
  wire[32:0] Switch_28_io_outPort_7;
  wire[32:0] Switch_28_io_outPort_6;
  wire[32:0] Switch_28_io_outPort_5;
  wire[32:0] Switch_28_io_outPort_4;
  wire[32:0] Switch_28_io_outPort_3;
  wire[32:0] Switch_28_io_outPort_2;
  wire[32:0] Switch_28_io_outPort_1;
  wire[32:0] Switch_28_io_outPort_0;
  wire[7:0] Switch_28_io_deqValid;
  wire[7:0] Switch_28_io_enqRdy;
  wire[23:0] Switch_28_io_outCUConfig;
  wire Switch_28_io_enqOR;
  wire[32:0] Switch_29_io_outPort_7;
  wire[32:0] Switch_29_io_outPort_6;
  wire[32:0] Switch_29_io_outPort_3;
  wire[32:0] Switch_29_io_outPort_2;
  wire[32:0] Switch_29_io_outPort_1;
  wire[32:0] Switch_29_io_outPort_0;
  wire[7:0] Switch_29_io_deqValid;
  wire[7:0] Switch_29_io_enqRdy;
  wire Switch_29_io_enqOR;
  wire[32:0] Switch_30_io_outPort_5;
  wire[32:0] Switch_30_io_outPort_3;
  wire[32:0] Switch_30_io_outPort_2;
  wire[32:0] Switch_30_io_outPort_1;
  wire[7:0] Switch_30_io_deqValid;
  wire[7:0] Switch_30_io_enqRdy;
  wire[32:0] Switch_31_io_outPort_6;
  wire[32:0] Switch_31_io_outPort_5;
  wire[32:0] Switch_31_io_outPort_3;
  wire[32:0] Switch_31_io_outPort_2;
  wire[32:0] Switch_31_io_outPort_1;
  wire[32:0] Switch_31_io_outPort_0;
  wire[7:0] Switch_31_io_deqValid;
  wire[7:0] Switch_31_io_enqRdy;
  wire Switch_31_io_enqOR;
  wire[32:0] Switch_32_io_outPort_6;
  wire[32:0] Switch_32_io_outPort_5;
  wire[32:0] Switch_32_io_outPort_3;
  wire[32:0] Switch_32_io_outPort_2;
  wire[32:0] Switch_32_io_outPort_1;
  wire[32:0] Switch_32_io_outPort_0;
  wire[7:0] Switch_32_io_deqValid;
  wire[7:0] Switch_32_io_enqRdy;
  wire Switch_32_io_enqOR;
  wire[32:0] Switch_33_io_outPort_6;
  wire[32:0] Switch_33_io_outPort_5;
  wire[32:0] Switch_33_io_outPort_3;
  wire[32:0] Switch_33_io_outPort_2;
  wire[32:0] Switch_33_io_outPort_1;
  wire[32:0] Switch_33_io_outPort_0;
  wire[7:0] Switch_33_io_deqValid;
  wire[7:0] Switch_33_io_enqRdy;
  wire Switch_33_io_enqOR;
  wire[32:0] Switch_34_io_outPort_6;
  wire[32:0] Switch_34_io_outPort_5;
  wire[32:0] Switch_34_io_outPort_3;
  wire[32:0] Switch_34_io_outPort_2;
  wire[32:0] Switch_34_io_outPort_1;
  wire[32:0] Switch_34_io_outPort_0;
  wire[7:0] Switch_34_io_deqValid;
  wire[7:0] Switch_34_io_enqRdy;
  wire Switch_34_io_enqOR;
  wire[32:0] Switch_35_io_outPort_6;
  wire[32:0] Switch_35_io_outPort_3;
  wire[32:0] Switch_35_io_outPort_2;
  wire[32:0] Switch_35_io_outPort_1;
  wire[7:0] Switch_35_io_deqValid;
  wire[7:0] Switch_35_io_enqRdy;
  wire Switch_35_io_enqOR;


  assign T0 = {1'h1, T1};
  assign T1 = {CU_24_io_enqRdyOut, 2'h3};
  assign T2 = {T8, T3};
  assign T3 = {T5, T4};
  assign T4 = {io_deqValid_10, 1'h0};
  assign T5 = {T7, T6};
  assign T6 = Switch_29_io_deqValid[1'h0:1'h0];
  assign T7 = Switch_34_io_deqValid[1'h1:1'h1];
  assign T8 = {1'h0, T9};
  assign T9 = {CU_24_io_deqValid, 2'h0};
  assign T10 = {T16, T11};
  assign T11 = {T13, T12};
  assign T12 = {io_enqRdy_10, 1'h1};
  assign T13 = {T15, T14};
  assign T14 = Switch_29_io_enqRdy[1'h0:1'h0];
  assign T15 = Switch_34_io_enqRdy[1'h1:1'h1];
  assign T16 = {1'h1, T17};
  assign T17 = {CU_24_io_enqRdy, 2'h3};
  assign T18 = {T20, T19};
  assign T19 = {CU_24_io_enqRdyOut, 1'h1};
  assign T20 = {1'h1, CU_23_io_enqRdyOut};
  assign T21 = {T28, T22};
  assign T22 = {T25, T23};
  assign T23 = {T24, io_deqValid_9};
  assign T24 = Switch_35_io_deqValid[2'h3:2'h3];
  assign T25 = {T27, T26};
  assign T26 = Switch_28_io_deqValid[1'h0:1'h0];
  assign T27 = Switch_33_io_deqValid[1'h1:1'h1];
  assign T28 = {T30, T29};
  assign T29 = {CU_24_io_deqValid, 1'h0};
  assign T30 = {1'h0, CU_23_io_deqValid};
  assign T31 = {T38, T32};
  assign T32 = {T35, T33};
  assign T33 = {T34, io_enqRdy_9};
  assign T34 = Switch_35_io_enqRdy[2'h3:2'h3];
  assign T35 = {T37, T36};
  assign T36 = Switch_28_io_enqRdy[1'h0:1'h0];
  assign T37 = Switch_33_io_enqRdy[1'h1:1'h1];
  assign T38 = {T40, T39};
  assign T39 = {CU_24_io_enqRdy, 1'h1};
  assign T40 = {1'h1, CU_23_io_enqRdy};
  assign T41 = {T43, T42};
  assign T42 = {CU_23_io_enqRdyOut, 1'h1};
  assign T43 = {1'h1, CU_22_io_enqRdyOut};
  assign T44 = {T51, T45};
  assign T45 = {T48, T46};
  assign T46 = {T47, io_deqValid_8};
  assign T47 = Switch_34_io_deqValid[2'h3:2'h3];
  assign T48 = {T50, T49};
  assign T49 = Switch_27_io_deqValid[1'h0:1'h0];
  assign T50 = Switch_32_io_deqValid[1'h1:1'h1];
  assign T51 = {T53, T52};
  assign T52 = {CU_23_io_deqValid, 1'h0};
  assign T53 = {1'h0, CU_22_io_deqValid};
  assign T54 = {T61, T55};
  assign T55 = {T58, T56};
  assign T56 = {T57, io_enqRdy_8};
  assign T57 = Switch_34_io_enqRdy[2'h3:2'h3];
  assign T58 = {T60, T59};
  assign T59 = Switch_27_io_enqRdy[1'h0:1'h0];
  assign T60 = Switch_32_io_enqRdy[1'h1:1'h1];
  assign T61 = {T63, T62};
  assign T62 = {CU_23_io_enqRdy, 1'h1};
  assign T63 = {1'h1, CU_22_io_enqRdy};
  assign T64 = {T66, T65};
  assign T65 = {CU_22_io_enqRdyOut, 1'h1};
  assign T66 = {1'h1, CU_21_io_enqRdyOut};
  assign T67 = {T74, T68};
  assign T68 = {T71, T69};
  assign T69 = {T70, io_deqValid_7};
  assign T70 = Switch_33_io_deqValid[2'h3:2'h3];
  assign T71 = {T73, T72};
  assign T72 = Switch_26_io_deqValid[1'h0:1'h0];
  assign T73 = Switch_31_io_deqValid[1'h1:1'h1];
  assign T74 = {T76, T75};
  assign T75 = {CU_22_io_deqValid, 1'h0};
  assign T76 = {1'h0, CU_21_io_deqValid};
  assign T77 = {T84, T78};
  assign T78 = {T81, T79};
  assign T79 = {T80, io_enqRdy_7};
  assign T80 = Switch_33_io_enqRdy[2'h3:2'h3];
  assign T81 = {T83, T82};
  assign T82 = Switch_26_io_enqRdy[1'h0:1'h0];
  assign T83 = Switch_31_io_enqRdy[1'h1:1'h1];
  assign T84 = {T86, T85};
  assign T85 = {CU_22_io_enqRdy, 1'h1};
  assign T86 = {1'h1, CU_21_io_enqRdy};
  assign T87 = {T89, T88};
  assign T88 = {CU_21_io_enqRdyOut, 1'h1};
  assign T89 = {1'h1, CU_20_io_enqRdyOut};
  assign T90 = {T97, T91};
  assign T91 = {T94, T92};
  assign T92 = {T93, io_deqValid_6};
  assign T93 = Switch_32_io_deqValid[2'h3:2'h3];
  assign T94 = {T96, T95};
  assign T95 = Switch_25_io_deqValid[1'h0:1'h0];
  assign T96 = Switch_30_io_deqValid[1'h1:1'h1];
  assign T97 = {T99, T98};
  assign T98 = {CU_21_io_deqValid, 1'h0};
  assign T99 = {1'h0, CU_20_io_deqValid};
  assign T100 = {T107, T101};
  assign T101 = {T104, T102};
  assign T102 = {T103, io_enqRdy_6};
  assign T103 = Switch_32_io_enqRdy[2'h3:2'h3];
  assign T104 = {T106, T105};
  assign T105 = Switch_25_io_enqRdy[1'h0:1'h0];
  assign T106 = Switch_30_io_enqRdy[1'h1:1'h1];
  assign T107 = {T109, T108};
  assign T108 = {CU_21_io_enqRdy, 1'h1};
  assign T109 = {1'h1, CU_20_io_enqRdy};
  assign T110 = {2'h3, T111};
  assign T111 = {CU_20_io_enqRdyOut, 1'h1};
  assign T112 = {T118, T113};
  assign T113 = {T116, T114};
  assign T114 = {T115, 1'h0};
  assign T115 = Switch_31_io_deqValid[2'h3:2'h3];
  assign T116 = {io_deqValid_5, T117};
  assign T117 = Switch_24_io_deqValid[1'h0:1'h0];
  assign T118 = {2'h0, T119};
  assign T119 = {CU_20_io_deqValid, 1'h0};
  assign T120 = {T126, T121};
  assign T121 = {T124, T122};
  assign T122 = {T123, 1'h1};
  assign T123 = Switch_31_io_enqRdy[2'h3:2'h3];
  assign T124 = {io_enqRdy_5, T125};
  assign T125 = Switch_24_io_enqRdy[1'h0:1'h0];
  assign T126 = {2'h3, T127};
  assign T127 = {CU_20_io_enqRdy, 1'h1};
  assign T128 = {CU_24_io_enqRdyOut, T129};
  assign T129 = {CU_19_io_enqRdyOut, 2'h3};
  assign T130 = {T137, T131};
  assign T131 = {T134, T132};
  assign T132 = {io_deqValid_11, T133};
  assign T133 = Switch_35_io_deqValid[2'h2:2'h2];
  assign T134 = {T136, T135};
  assign T135 = Switch_23_io_deqValid[1'h0:1'h0];
  assign T136 = Switch_28_io_deqValid[1'h1:1'h1];
  assign T137 = {CU_24_io_deqValid, T138};
  assign T138 = {CU_19_io_deqValid, 2'h0};
  assign T139 = {T146, T140};
  assign T140 = {T143, T141};
  assign T141 = {io_enqRdy_11, T142};
  assign T142 = Switch_35_io_enqRdy[2'h2:2'h2];
  assign T143 = {T145, T144};
  assign T144 = Switch_23_io_enqRdy[1'h0:1'h0];
  assign T145 = Switch_28_io_enqRdy[1'h1:1'h1];
  assign T146 = {CU_24_io_enqRdy, T147};
  assign T147 = {CU_19_io_enqRdy, 2'h3};
  assign T148 = {T150, T149};
  assign T149 = {CU_19_io_enqRdyOut, CU_24_io_enqRdyOut};
  assign T150 = {CU_23_io_enqRdyOut, CU_18_io_enqRdyOut};
  assign T151 = {T159, T152};
  assign T152 = {T156, T153};
  assign T153 = {T155, T154};
  assign T154 = Switch_34_io_deqValid[2'h2:2'h2];
  assign T155 = Switch_29_io_deqValid[2'h3:2'h3];
  assign T156 = {T158, T157};
  assign T157 = Switch_22_io_deqValid[1'h0:1'h0];
  assign T158 = Switch_27_io_deqValid[1'h1:1'h1];
  assign T159 = {T161, T160};
  assign T160 = {CU_19_io_deqValid, CU_24_io_deqValid};
  assign T161 = {CU_23_io_deqValid, CU_18_io_deqValid};
  assign T162 = {T170, T163};
  assign T163 = {T167, T164};
  assign T164 = {T166, T165};
  assign T165 = Switch_34_io_enqRdy[2'h2:2'h2];
  assign T166 = Switch_29_io_enqRdy[2'h3:2'h3];
  assign T167 = {T169, T168};
  assign T168 = Switch_22_io_enqRdy[1'h0:1'h0];
  assign T169 = Switch_27_io_enqRdy[1'h1:1'h1];
  assign T170 = {T172, T171};
  assign T171 = {CU_19_io_enqRdy, CU_24_io_enqRdy};
  assign T172 = {CU_23_io_enqRdy, CU_18_io_enqRdy};
  assign T173 = {T175, T174};
  assign T174 = {CU_18_io_enqRdyOut, CU_23_io_enqRdyOut};
  assign T175 = {CU_22_io_enqRdyOut, CU_17_io_enqRdyOut};
  assign T176 = {T184, T177};
  assign T177 = {T181, T178};
  assign T178 = {T180, T179};
  assign T179 = Switch_33_io_deqValid[2'h2:2'h2];
  assign T180 = Switch_28_io_deqValid[2'h3:2'h3];
  assign T181 = {T183, T182};
  assign T182 = Switch_21_io_deqValid[1'h0:1'h0];
  assign T183 = Switch_26_io_deqValid[1'h1:1'h1];
  assign T184 = {T186, T185};
  assign T185 = {CU_18_io_deqValid, CU_23_io_deqValid};
  assign T186 = {CU_22_io_deqValid, CU_17_io_deqValid};
  assign T187 = {T195, T188};
  assign T188 = {T192, T189};
  assign T189 = {T191, T190};
  assign T190 = Switch_33_io_enqRdy[2'h2:2'h2];
  assign T191 = Switch_28_io_enqRdy[2'h3:2'h3];
  assign T192 = {T194, T193};
  assign T193 = Switch_21_io_enqRdy[1'h0:1'h0];
  assign T194 = Switch_26_io_enqRdy[1'h1:1'h1];
  assign T195 = {T197, T196};
  assign T196 = {CU_18_io_enqRdy, CU_23_io_enqRdy};
  assign T197 = {CU_22_io_enqRdy, CU_17_io_enqRdy};
  assign T198 = {T200, T199};
  assign T199 = {CU_17_io_enqRdyOut, CU_22_io_enqRdyOut};
  assign T200 = {CU_21_io_enqRdyOut, CU_16_io_enqRdyOut};
  assign T201 = {T209, T202};
  assign T202 = {T206, T203};
  assign T203 = {T205, T204};
  assign T204 = Switch_32_io_deqValid[2'h2:2'h2];
  assign T205 = Switch_27_io_deqValid[2'h3:2'h3];
  assign T206 = {T208, T207};
  assign T207 = Switch_20_io_deqValid[1'h0:1'h0];
  assign T208 = Switch_25_io_deqValid[1'h1:1'h1];
  assign T209 = {T211, T210};
  assign T210 = {CU_17_io_deqValid, CU_22_io_deqValid};
  assign T211 = {CU_21_io_deqValid, CU_16_io_deqValid};
  assign T212 = {T220, T213};
  assign T213 = {T217, T214};
  assign T214 = {T216, T215};
  assign T215 = Switch_32_io_enqRdy[2'h2:2'h2];
  assign T216 = Switch_27_io_enqRdy[2'h3:2'h3];
  assign T217 = {T219, T218};
  assign T218 = Switch_20_io_enqRdy[1'h0:1'h0];
  assign T219 = Switch_25_io_enqRdy[1'h1:1'h1];
  assign T220 = {T222, T221};
  assign T221 = {CU_17_io_enqRdy, CU_22_io_enqRdy};
  assign T222 = {CU_21_io_enqRdy, CU_16_io_enqRdy};
  assign T223 = {T225, T224};
  assign T224 = {CU_16_io_enqRdyOut, CU_21_io_enqRdyOut};
  assign T225 = {CU_20_io_enqRdyOut, CU_15_io_enqRdyOut};
  assign T226 = {T234, T227};
  assign T227 = {T231, T228};
  assign T228 = {T230, T229};
  assign T229 = Switch_31_io_deqValid[2'h2:2'h2];
  assign T230 = Switch_26_io_deqValid[2'h3:2'h3];
  assign T231 = {T233, T232};
  assign T232 = Switch_19_io_deqValid[1'h0:1'h0];
  assign T233 = Switch_24_io_deqValid[1'h1:1'h1];
  assign T234 = {T236, T235};
  assign T235 = {CU_16_io_deqValid, CU_21_io_deqValid};
  assign T236 = {CU_20_io_deqValid, CU_15_io_deqValid};
  assign T237 = {T245, T238};
  assign T238 = {T242, T239};
  assign T239 = {T241, T240};
  assign T240 = Switch_31_io_enqRdy[2'h2:2'h2];
  assign T241 = Switch_26_io_enqRdy[2'h3:2'h3];
  assign T242 = {T244, T243};
  assign T243 = Switch_19_io_enqRdy[1'h0:1'h0];
  assign T244 = Switch_24_io_enqRdy[1'h1:1'h1];
  assign T245 = {T247, T246};
  assign T246 = {CU_16_io_enqRdy, CU_21_io_enqRdy};
  assign T247 = {CU_20_io_enqRdy, CU_15_io_enqRdy};
  assign T248 = {2'h3, T249};
  assign T249 = {CU_15_io_enqRdyOut, CU_20_io_enqRdyOut};
  assign T250 = {T257, T251};
  assign T251 = {T255, T252};
  assign T252 = {T254, T253};
  assign T253 = Switch_30_io_deqValid[2'h2:2'h2];
  assign T254 = Switch_25_io_deqValid[2'h3:2'h3];
  assign T255 = {io_deqValid_4, T256};
  assign T256 = Switch_18_io_deqValid[1'h0:1'h0];
  assign T257 = {2'h0, T258};
  assign T258 = {CU_15_io_deqValid, CU_20_io_deqValid};
  assign T259 = {T266, T260};
  assign T260 = {T264, T261};
  assign T261 = {T263, T262};
  assign T262 = Switch_30_io_enqRdy[2'h2:2'h2];
  assign T263 = Switch_25_io_enqRdy[2'h3:2'h3];
  assign T264 = {io_enqRdy_4, T265};
  assign T265 = Switch_18_io_enqRdy[1'h0:1'h0];
  assign T266 = {2'h3, T267};
  assign T267 = {CU_15_io_enqRdy, CU_20_io_enqRdy};
  assign T268 = {CU_19_io_enqRdyOut, T269};
  assign T269 = {CU_14_io_enqRdyOut, 2'h3};
  assign T270 = {T277, T271};
  assign T271 = {T274, T272};
  assign T272 = {io_deqValid_12, T273};
  assign T273 = Switch_29_io_deqValid[2'h2:2'h2];
  assign T274 = {T276, T275};
  assign T275 = Switch_17_io_deqValid[1'h0:1'h0];
  assign T276 = Switch_22_io_deqValid[1'h1:1'h1];
  assign T277 = {CU_19_io_deqValid, T278};
  assign T278 = {CU_14_io_deqValid, 2'h0};
  assign T279 = {T286, T280};
  assign T280 = {T283, T281};
  assign T281 = {io_enqRdy_12, T282};
  assign T282 = Switch_29_io_enqRdy[2'h2:2'h2];
  assign T283 = {T285, T284};
  assign T284 = Switch_17_io_enqRdy[1'h0:1'h0];
  assign T285 = Switch_22_io_enqRdy[1'h1:1'h1];
  assign T286 = {CU_19_io_enqRdy, T287};
  assign T287 = {CU_14_io_enqRdy, 2'h3};
  assign T288 = {T290, T289};
  assign T289 = {CU_14_io_enqRdyOut, CU_19_io_enqRdyOut};
  assign T290 = {CU_18_io_enqRdyOut, CU_13_io_enqRdyOut};
  assign T291 = {T299, T292};
  assign T292 = {T296, T293};
  assign T293 = {T295, T294};
  assign T294 = Switch_28_io_deqValid[2'h2:2'h2];
  assign T295 = Switch_23_io_deqValid[2'h3:2'h3];
  assign T296 = {T298, T297};
  assign T297 = Switch_16_io_deqValid[1'h0:1'h0];
  assign T298 = Switch_21_io_deqValid[1'h1:1'h1];
  assign T299 = {T301, T300};
  assign T300 = {CU_14_io_deqValid, CU_19_io_deqValid};
  assign T301 = {CU_18_io_deqValid, CU_13_io_deqValid};
  assign T302 = {T310, T303};
  assign T303 = {T307, T304};
  assign T304 = {T306, T305};
  assign T305 = Switch_28_io_enqRdy[2'h2:2'h2];
  assign T306 = Switch_23_io_enqRdy[2'h3:2'h3];
  assign T307 = {T309, T308};
  assign T308 = Switch_16_io_enqRdy[1'h0:1'h0];
  assign T309 = Switch_21_io_enqRdy[1'h1:1'h1];
  assign T310 = {T312, T311};
  assign T311 = {CU_14_io_enqRdy, CU_19_io_enqRdy};
  assign T312 = {CU_18_io_enqRdy, CU_13_io_enqRdy};
  assign T313 = {T315, T314};
  assign T314 = {CU_13_io_enqRdyOut, CU_18_io_enqRdyOut};
  assign T315 = {CU_17_io_enqRdyOut, CU_12_io_enqRdyOut};
  assign T316 = {T324, T317};
  assign T317 = {T321, T318};
  assign T318 = {T320, T319};
  assign T319 = Switch_27_io_deqValid[2'h2:2'h2];
  assign T320 = Switch_22_io_deqValid[2'h3:2'h3];
  assign T321 = {T323, T322};
  assign T322 = Switch_15_io_deqValid[1'h0:1'h0];
  assign T323 = Switch_20_io_deqValid[1'h1:1'h1];
  assign T324 = {T326, T325};
  assign T325 = {CU_13_io_deqValid, CU_18_io_deqValid};
  assign T326 = {CU_17_io_deqValid, CU_12_io_deqValid};
  assign T327 = {T335, T328};
  assign T328 = {T332, T329};
  assign T329 = {T331, T330};
  assign T330 = Switch_27_io_enqRdy[2'h2:2'h2];
  assign T331 = Switch_22_io_enqRdy[2'h3:2'h3];
  assign T332 = {T334, T333};
  assign T333 = Switch_15_io_enqRdy[1'h0:1'h0];
  assign T334 = Switch_20_io_enqRdy[1'h1:1'h1];
  assign T335 = {T337, T336};
  assign T336 = {CU_13_io_enqRdy, CU_18_io_enqRdy};
  assign T337 = {CU_17_io_enqRdy, CU_12_io_enqRdy};
  assign T338 = {T340, T339};
  assign T339 = {CU_12_io_enqRdyOut, CU_17_io_enqRdyOut};
  assign T340 = {CU_16_io_enqRdyOut, CU_11_io_enqRdyOut};
  assign T341 = {T349, T342};
  assign T342 = {T346, T343};
  assign T343 = {T345, T344};
  assign T344 = Switch_26_io_deqValid[2'h2:2'h2];
  assign T345 = Switch_21_io_deqValid[2'h3:2'h3];
  assign T346 = {T348, T347};
  assign T347 = Switch_14_io_deqValid[1'h0:1'h0];
  assign T348 = Switch_19_io_deqValid[1'h1:1'h1];
  assign T349 = {T351, T350};
  assign T350 = {CU_12_io_deqValid, CU_17_io_deqValid};
  assign T351 = {CU_16_io_deqValid, CU_11_io_deqValid};
  assign T352 = {T360, T353};
  assign T353 = {T357, T354};
  assign T354 = {T356, T355};
  assign T355 = Switch_26_io_enqRdy[2'h2:2'h2];
  assign T356 = Switch_21_io_enqRdy[2'h3:2'h3];
  assign T357 = {T359, T358};
  assign T358 = Switch_14_io_enqRdy[1'h0:1'h0];
  assign T359 = Switch_19_io_enqRdy[1'h1:1'h1];
  assign T360 = {T362, T361};
  assign T361 = {CU_12_io_enqRdy, CU_17_io_enqRdy};
  assign T362 = {CU_16_io_enqRdy, CU_11_io_enqRdy};
  assign T363 = {T365, T364};
  assign T364 = {CU_11_io_enqRdyOut, CU_16_io_enqRdyOut};
  assign T365 = {CU_15_io_enqRdyOut, CU_10_io_enqRdyOut};
  assign T366 = {T374, T367};
  assign T367 = {T371, T368};
  assign T368 = {T370, T369};
  assign T369 = Switch_25_io_deqValid[2'h2:2'h2];
  assign T370 = Switch_20_io_deqValid[2'h3:2'h3];
  assign T371 = {T373, T372};
  assign T372 = Switch_13_io_deqValid[1'h0:1'h0];
  assign T373 = Switch_18_io_deqValid[1'h1:1'h1];
  assign T374 = {T376, T375};
  assign T375 = {CU_11_io_deqValid, CU_16_io_deqValid};
  assign T376 = {CU_15_io_deqValid, CU_10_io_deqValid};
  assign T377 = {T385, T378};
  assign T378 = {T382, T379};
  assign T379 = {T381, T380};
  assign T380 = Switch_25_io_enqRdy[2'h2:2'h2];
  assign T381 = Switch_20_io_enqRdy[2'h3:2'h3];
  assign T382 = {T384, T383};
  assign T383 = Switch_13_io_enqRdy[1'h0:1'h0];
  assign T384 = Switch_18_io_enqRdy[1'h1:1'h1];
  assign T385 = {T387, T386};
  assign T386 = {CU_11_io_enqRdy, CU_16_io_enqRdy};
  assign T387 = {CU_15_io_enqRdy, CU_10_io_enqRdy};
  assign T388 = {2'h3, T389};
  assign T389 = {CU_10_io_enqRdyOut, CU_15_io_enqRdyOut};
  assign T390 = {T397, T391};
  assign T391 = {T395, T392};
  assign T392 = {T394, T393};
  assign T393 = Switch_24_io_deqValid[2'h2:2'h2];
  assign T394 = Switch_19_io_deqValid[2'h3:2'h3];
  assign T395 = {io_deqValid_3, T396};
  assign T396 = Switch_12_io_deqValid[1'h0:1'h0];
  assign T397 = {2'h0, T398};
  assign T398 = {CU_10_io_deqValid, CU_15_io_deqValid};
  assign T399 = {T406, T400};
  assign T400 = {T404, T401};
  assign T401 = {T403, T402};
  assign T402 = Switch_24_io_enqRdy[2'h2:2'h2];
  assign T403 = Switch_19_io_enqRdy[2'h3:2'h3];
  assign T404 = {io_enqRdy_3, T405};
  assign T405 = Switch_12_io_enqRdy[1'h0:1'h0];
  assign T406 = {2'h3, T407};
  assign T407 = {CU_10_io_enqRdy, CU_15_io_enqRdy};
  assign T408 = {CU_14_io_enqRdyOut, T409};
  assign T409 = {CU_9_io_enqRdyOut, 2'h3};
  assign T410 = {T417, T411};
  assign T411 = {T414, T412};
  assign T412 = {io_deqValid_13, T413};
  assign T413 = Switch_23_io_deqValid[2'h2:2'h2];
  assign T414 = {T416, T415};
  assign T415 = Switch_11_io_deqValid[1'h0:1'h0];
  assign T416 = Switch_16_io_deqValid[1'h1:1'h1];
  assign T417 = {CU_14_io_deqValid, T418};
  assign T418 = {CU_9_io_deqValid, 2'h0};
  assign T419 = {T426, T420};
  assign T420 = {T423, T421};
  assign T421 = {io_enqRdy_13, T422};
  assign T422 = Switch_23_io_enqRdy[2'h2:2'h2];
  assign T423 = {T425, T424};
  assign T424 = Switch_11_io_enqRdy[1'h0:1'h0];
  assign T425 = Switch_16_io_enqRdy[1'h1:1'h1];
  assign T426 = {CU_14_io_enqRdy, T427};
  assign T427 = {CU_9_io_enqRdy, 2'h3};
  assign T428 = {T430, T429};
  assign T429 = {CU_9_io_enqRdyOut, CU_14_io_enqRdyOut};
  assign T430 = {CU_13_io_enqRdyOut, CU_8_io_enqRdyOut};
  assign T431 = {T439, T432};
  assign T432 = {T436, T433};
  assign T433 = {T435, T434};
  assign T434 = Switch_22_io_deqValid[2'h2:2'h2];
  assign T435 = Switch_17_io_deqValid[2'h3:2'h3];
  assign T436 = {T438, T437};
  assign T437 = Switch_10_io_deqValid[1'h0:1'h0];
  assign T438 = Switch_15_io_deqValid[1'h1:1'h1];
  assign T439 = {T441, T440};
  assign T440 = {CU_9_io_deqValid, CU_14_io_deqValid};
  assign T441 = {CU_13_io_deqValid, CU_8_io_deqValid};
  assign T442 = {T450, T443};
  assign T443 = {T447, T444};
  assign T444 = {T446, T445};
  assign T445 = Switch_22_io_enqRdy[2'h2:2'h2];
  assign T446 = Switch_17_io_enqRdy[2'h3:2'h3];
  assign T447 = {T449, T448};
  assign T448 = Switch_10_io_enqRdy[1'h0:1'h0];
  assign T449 = Switch_15_io_enqRdy[1'h1:1'h1];
  assign T450 = {T452, T451};
  assign T451 = {CU_9_io_enqRdy, CU_14_io_enqRdy};
  assign T452 = {CU_13_io_enqRdy, CU_8_io_enqRdy};
  assign T453 = {T455, T454};
  assign T454 = {CU_8_io_enqRdyOut, CU_13_io_enqRdyOut};
  assign T455 = {CU_12_io_enqRdyOut, CU_7_io_enqRdyOut};
  assign T456 = {T464, T457};
  assign T457 = {T461, T458};
  assign T458 = {T460, T459};
  assign T459 = Switch_21_io_deqValid[2'h2:2'h2];
  assign T460 = Switch_16_io_deqValid[2'h3:2'h3];
  assign T461 = {T463, T462};
  assign T462 = Switch_9_io_deqValid[1'h0:1'h0];
  assign T463 = Switch_14_io_deqValid[1'h1:1'h1];
  assign T464 = {T466, T465};
  assign T465 = {CU_8_io_deqValid, CU_13_io_deqValid};
  assign T466 = {CU_12_io_deqValid, CU_7_io_deqValid};
  assign T467 = {T475, T468};
  assign T468 = {T472, T469};
  assign T469 = {T471, T470};
  assign T470 = Switch_21_io_enqRdy[2'h2:2'h2];
  assign T471 = Switch_16_io_enqRdy[2'h3:2'h3];
  assign T472 = {T474, T473};
  assign T473 = Switch_9_io_enqRdy[1'h0:1'h0];
  assign T474 = Switch_14_io_enqRdy[1'h1:1'h1];
  assign T475 = {T477, T476};
  assign T476 = {CU_8_io_enqRdy, CU_13_io_enqRdy};
  assign T477 = {CU_12_io_enqRdy, CU_7_io_enqRdy};
  assign T478 = {T480, T479};
  assign T479 = {CU_7_io_enqRdyOut, CU_12_io_enqRdyOut};
  assign T480 = {CU_11_io_enqRdyOut, CU_6_io_enqRdyOut};
  assign T481 = {T489, T482};
  assign T482 = {T486, T483};
  assign T483 = {T485, T484};
  assign T484 = Switch_20_io_deqValid[2'h2:2'h2];
  assign T485 = Switch_15_io_deqValid[2'h3:2'h3];
  assign T486 = {T488, T487};
  assign T487 = Switch_8_io_deqValid[1'h0:1'h0];
  assign T488 = Switch_13_io_deqValid[1'h1:1'h1];
  assign T489 = {T491, T490};
  assign T490 = {CU_7_io_deqValid, CU_12_io_deqValid};
  assign T491 = {CU_11_io_deqValid, CU_6_io_deqValid};
  assign T492 = {T500, T493};
  assign T493 = {T497, T494};
  assign T494 = {T496, T495};
  assign T495 = Switch_20_io_enqRdy[2'h2:2'h2];
  assign T496 = Switch_15_io_enqRdy[2'h3:2'h3];
  assign T497 = {T499, T498};
  assign T498 = Switch_8_io_enqRdy[1'h0:1'h0];
  assign T499 = Switch_13_io_enqRdy[1'h1:1'h1];
  assign T500 = {T502, T501};
  assign T501 = {CU_7_io_enqRdy, CU_12_io_enqRdy};
  assign T502 = {CU_11_io_enqRdy, CU_6_io_enqRdy};
  assign T503 = {T505, T504};
  assign T504 = {CU_6_io_enqRdyOut, CU_11_io_enqRdyOut};
  assign T505 = {CU_10_io_enqRdyOut, CU_5_io_enqRdyOut};
  assign T506 = {T514, T507};
  assign T507 = {T511, T508};
  assign T508 = {T510, T509};
  assign T509 = Switch_19_io_deqValid[2'h2:2'h2];
  assign T510 = Switch_14_io_deqValid[2'h3:2'h3];
  assign T511 = {T513, T512};
  assign T512 = Switch_7_io_deqValid[1'h0:1'h0];
  assign T513 = Switch_12_io_deqValid[1'h1:1'h1];
  assign T514 = {T516, T515};
  assign T515 = {CU_6_io_deqValid, CU_11_io_deqValid};
  assign T516 = {CU_10_io_deqValid, CU_5_io_deqValid};
  assign T517 = {T525, T518};
  assign T518 = {T522, T519};
  assign T519 = {T521, T520};
  assign T520 = Switch_19_io_enqRdy[2'h2:2'h2];
  assign T521 = Switch_14_io_enqRdy[2'h3:2'h3];
  assign T522 = {T524, T523};
  assign T523 = Switch_7_io_enqRdy[1'h0:1'h0];
  assign T524 = Switch_12_io_enqRdy[1'h1:1'h1];
  assign T525 = {T527, T526};
  assign T526 = {CU_6_io_enqRdy, CU_11_io_enqRdy};
  assign T527 = {CU_10_io_enqRdy, CU_5_io_enqRdy};
  assign T528 = {2'h3, T529};
  assign T529 = {CU_5_io_enqRdyOut, CU_10_io_enqRdyOut};
  assign T530 = {T537, T531};
  assign T531 = {T535, T532};
  assign T532 = {T534, T533};
  assign T533 = Switch_18_io_deqValid[2'h2:2'h2];
  assign T534 = Switch_13_io_deqValid[2'h3:2'h3];
  assign T535 = {io_deqValid_2, T536};
  assign T536 = Switch_6_io_deqValid[1'h0:1'h0];
  assign T537 = {2'h0, T538};
  assign T538 = {CU_5_io_deqValid, CU_10_io_deqValid};
  assign T539 = {T546, T540};
  assign T540 = {T544, T541};
  assign T541 = {T543, T542};
  assign T542 = Switch_18_io_enqRdy[2'h2:2'h2];
  assign T543 = Switch_13_io_enqRdy[2'h3:2'h3];
  assign T544 = {io_enqRdy_2, T545};
  assign T545 = Switch_6_io_enqRdy[1'h0:1'h0];
  assign T546 = {2'h3, T547};
  assign T547 = {CU_5_io_enqRdy, CU_10_io_enqRdy};
  assign T548 = {CU_9_io_enqRdyOut, T549};
  assign T549 = {CU_4_io_enqRdyOut, 2'h3};
  assign T550 = {T557, T551};
  assign T551 = {T554, T552};
  assign T552 = {io_deqValid_14, T553};
  assign T553 = Switch_17_io_deqValid[2'h2:2'h2];
  assign T554 = {T556, T555};
  assign T555 = Switch_5_io_deqValid[1'h0:1'h0];
  assign T556 = Switch_10_io_deqValid[1'h1:1'h1];
  assign T557 = {CU_9_io_deqValid, T558};
  assign T558 = {CU_4_io_deqValid, 2'h0};
  assign T559 = {T566, T560};
  assign T560 = {T563, T561};
  assign T561 = {io_enqRdy_14, T562};
  assign T562 = Switch_17_io_enqRdy[2'h2:2'h2];
  assign T563 = {T565, T564};
  assign T564 = Switch_5_io_enqRdy[1'h0:1'h0];
  assign T565 = Switch_10_io_enqRdy[1'h1:1'h1];
  assign T566 = {CU_9_io_enqRdy, T567};
  assign T567 = {CU_4_io_enqRdy, 2'h3};
  assign T568 = {T570, T569};
  assign T569 = {CU_4_io_enqRdyOut, CU_9_io_enqRdyOut};
  assign T570 = {CU_8_io_enqRdyOut, CU_3_io_enqRdyOut};
  assign T571 = {T579, T572};
  assign T572 = {T576, T573};
  assign T573 = {T575, T574};
  assign T574 = Switch_16_io_deqValid[2'h2:2'h2];
  assign T575 = Switch_11_io_deqValid[2'h3:2'h3];
  assign T576 = {T578, T577};
  assign T577 = Switch_4_io_deqValid[1'h0:1'h0];
  assign T578 = Switch_9_io_deqValid[1'h1:1'h1];
  assign T579 = {T581, T580};
  assign T580 = {CU_4_io_deqValid, CU_9_io_deqValid};
  assign T581 = {CU_8_io_deqValid, CU_3_io_deqValid};
  assign T582 = {T590, T583};
  assign T583 = {T587, T584};
  assign T584 = {T586, T585};
  assign T585 = Switch_16_io_enqRdy[2'h2:2'h2];
  assign T586 = Switch_11_io_enqRdy[2'h3:2'h3];
  assign T587 = {T589, T588};
  assign T588 = Switch_4_io_enqRdy[1'h0:1'h0];
  assign T589 = Switch_9_io_enqRdy[1'h1:1'h1];
  assign T590 = {T592, T591};
  assign T591 = {CU_4_io_enqRdy, CU_9_io_enqRdy};
  assign T592 = {CU_8_io_enqRdy, CU_3_io_enqRdy};
  assign T593 = {T595, T594};
  assign T594 = {CU_3_io_enqRdyOut, CU_8_io_enqRdyOut};
  assign T595 = {CU_7_io_enqRdyOut, CU_2_io_enqRdyOut};
  assign T596 = {T604, T597};
  assign T597 = {T601, T598};
  assign T598 = {T600, T599};
  assign T599 = Switch_15_io_deqValid[2'h2:2'h2];
  assign T600 = Switch_10_io_deqValid[2'h3:2'h3];
  assign T601 = {T603, T602};
  assign T602 = Switch_3_io_deqValid[1'h0:1'h0];
  assign T603 = Switch_8_io_deqValid[1'h1:1'h1];
  assign T604 = {T606, T605};
  assign T605 = {CU_3_io_deqValid, CU_8_io_deqValid};
  assign T606 = {CU_7_io_deqValid, CU_2_io_deqValid};
  assign T607 = {T615, T608};
  assign T608 = {T612, T609};
  assign T609 = {T611, T610};
  assign T610 = Switch_15_io_enqRdy[2'h2:2'h2];
  assign T611 = Switch_10_io_enqRdy[2'h3:2'h3];
  assign T612 = {T614, T613};
  assign T613 = Switch_3_io_enqRdy[1'h0:1'h0];
  assign T614 = Switch_8_io_enqRdy[1'h1:1'h1];
  assign T615 = {T617, T616};
  assign T616 = {CU_3_io_enqRdy, CU_8_io_enqRdy};
  assign T617 = {CU_7_io_enqRdy, CU_2_io_enqRdy};
  assign T618 = {T620, T619};
  assign T619 = {CU_2_io_enqRdyOut, CU_7_io_enqRdyOut};
  assign T620 = {CU_6_io_enqRdyOut, CU_1_io_enqRdyOut};
  assign T621 = {T629, T622};
  assign T622 = {T626, T623};
  assign T623 = {T625, T624};
  assign T624 = Switch_14_io_deqValid[2'h2:2'h2];
  assign T625 = Switch_9_io_deqValid[2'h3:2'h3];
  assign T626 = {T628, T627};
  assign T627 = Switch_2_io_deqValid[1'h0:1'h0];
  assign T628 = Switch_7_io_deqValid[1'h1:1'h1];
  assign T629 = {T631, T630};
  assign T630 = {CU_2_io_deqValid, CU_7_io_deqValid};
  assign T631 = {CU_6_io_deqValid, CU_1_io_deqValid};
  assign T632 = {T640, T633};
  assign T633 = {T637, T634};
  assign T634 = {T636, T635};
  assign T635 = Switch_14_io_enqRdy[2'h2:2'h2];
  assign T636 = Switch_9_io_enqRdy[2'h3:2'h3];
  assign T637 = {T639, T638};
  assign T638 = Switch_2_io_enqRdy[1'h0:1'h0];
  assign T639 = Switch_7_io_enqRdy[1'h1:1'h1];
  assign T640 = {T642, T641};
  assign T641 = {CU_2_io_enqRdy, CU_7_io_enqRdy};
  assign T642 = {CU_6_io_enqRdy, CU_1_io_enqRdy};
  assign T643 = {T645, T644};
  assign T644 = {CU_1_io_enqRdyOut, CU_6_io_enqRdyOut};
  assign T645 = {CU_5_io_enqRdyOut, CU_io_enqRdyOut};
  assign T646 = {T654, T647};
  assign T647 = {T651, T648};
  assign T648 = {T650, T649};
  assign T649 = Switch_13_io_deqValid[2'h2:2'h2];
  assign T650 = Switch_8_io_deqValid[2'h3:2'h3];
  assign T651 = {T653, T652};
  assign T652 = Switch_1_io_deqValid[1'h0:1'h0];
  assign T653 = Switch_6_io_deqValid[1'h1:1'h1];
  assign T654 = {T656, T655};
  assign T655 = {CU_1_io_deqValid, CU_6_io_deqValid};
  assign T656 = {CU_5_io_deqValid, CU_io_deqValid};
  assign T657 = {T665, T658};
  assign T658 = {T662, T659};
  assign T659 = {T661, T660};
  assign T660 = Switch_13_io_enqRdy[2'h2:2'h2];
  assign T661 = Switch_8_io_enqRdy[2'h3:2'h3];
  assign T662 = {T664, T663};
  assign T663 = Switch_1_io_enqRdy[1'h0:1'h0];
  assign T664 = Switch_6_io_enqRdy[1'h1:1'h1];
  assign T665 = {T667, T666};
  assign T666 = {CU_1_io_enqRdy, CU_6_io_enqRdy};
  assign T667 = {CU_5_io_enqRdy, CU_io_enqRdy};
  assign T668 = {2'h3, T669};
  assign T669 = {CU_io_enqRdyOut, CU_5_io_enqRdyOut};
  assign T670 = {T677, T671};
  assign T671 = {T675, T672};
  assign T672 = {T674, T673};
  assign T673 = Switch_12_io_deqValid[2'h2:2'h2];
  assign T674 = Switch_7_io_deqValid[2'h3:2'h3];
  assign T675 = {io_deqValid_1, T676};
  assign T676 = Switch_io_deqValid[1'h0:1'h0];
  assign T677 = {2'h0, T678};
  assign T678 = {CU_io_deqValid, CU_5_io_deqValid};
  assign T679 = {T686, T680};
  assign T680 = {T684, T681};
  assign T681 = {T683, T682};
  assign T682 = Switch_12_io_enqRdy[2'h2:2'h2];
  assign T683 = Switch_7_io_enqRdy[2'h3:2'h3];
  assign T684 = {io_enqRdy_1, T685};
  assign T685 = Switch_io_enqRdy[1'h0:1'h0];
  assign T686 = {2'h3, T687};
  assign T687 = {CU_io_enqRdy, CU_5_io_enqRdy};
  assign T688 = {CU_4_io_enqRdyOut, 3'h7};
  assign T689 = {T693, T690};
  assign T690 = {1'h0, T691};
  assign T691 = {io_deqValid_15, T692};
  assign T692 = Switch_11_io_deqValid[2'h2:2'h2];
  assign T693 = {CU_4_io_deqValid, T694};
  assign T694 = {3'h0, T695};
  assign T695 = Switch_4_io_deqValid[1'h1:1'h1];
  assign T696 = {T700, T697};
  assign T697 = {1'h1, T698};
  assign T698 = {io_enqRdy_15, T699};
  assign T699 = Switch_11_io_enqRdy[2'h2:2'h2];
  assign T700 = {CU_4_io_enqRdy, T701};
  assign T701 = {3'h7, T702};
  assign T702 = Switch_4_io_enqRdy[1'h1:1'h1];
  assign T703 = {CU_3_io_enqRdyOut, T704};
  assign T704 = {2'h3, CU_4_io_enqRdyOut};
  assign T705 = {T712, T706};
  assign T706 = {T710, T707};
  assign T707 = {T709, T708};
  assign T708 = Switch_10_io_deqValid[2'h2:2'h2];
  assign T709 = Switch_5_io_deqValid[2'h3:2'h3];
  assign T710 = {T711, io_deqValid_16};
  assign T711 = Switch_3_io_deqValid[1'h1:1'h1];
  assign T712 = {CU_3_io_deqValid, T713};
  assign T713 = {2'h0, CU_4_io_deqValid};
  assign T714 = {T721, T715};
  assign T715 = {T719, T716};
  assign T716 = {T718, T717};
  assign T717 = Switch_10_io_enqRdy[2'h2:2'h2];
  assign T718 = Switch_5_io_enqRdy[2'h3:2'h3];
  assign T719 = {T720, io_enqRdy_16};
  assign T720 = Switch_3_io_enqRdy[1'h1:1'h1];
  assign T721 = {CU_3_io_enqRdy, T722};
  assign T722 = {2'h3, CU_4_io_enqRdy};
  assign T723 = {CU_2_io_enqRdyOut, T724};
  assign T724 = {2'h3, CU_3_io_enqRdyOut};
  assign T725 = {T732, T726};
  assign T726 = {T730, T727};
  assign T727 = {T729, T728};
  assign T728 = Switch_9_io_deqValid[2'h2:2'h2];
  assign T729 = Switch_4_io_deqValid[2'h3:2'h3];
  assign T730 = {T731, io_deqValid_17};
  assign T731 = Switch_2_io_deqValid[1'h1:1'h1];
  assign T732 = {CU_2_io_deqValid, T733};
  assign T733 = {2'h0, CU_3_io_deqValid};
  assign T734 = {T741, T735};
  assign T735 = {T739, T736};
  assign T736 = {T738, T737};
  assign T737 = Switch_9_io_enqRdy[2'h2:2'h2];
  assign T738 = Switch_4_io_enqRdy[2'h3:2'h3];
  assign T739 = {T740, io_enqRdy_17};
  assign T740 = Switch_2_io_enqRdy[1'h1:1'h1];
  assign T741 = {CU_2_io_enqRdy, T742};
  assign T742 = {2'h3, CU_3_io_enqRdy};
  assign T743 = {CU_1_io_enqRdyOut, T744};
  assign T744 = {2'h3, CU_2_io_enqRdyOut};
  assign T745 = {T752, T746};
  assign T746 = {T750, T747};
  assign T747 = {T749, T748};
  assign T748 = Switch_8_io_deqValid[2'h2:2'h2];
  assign T749 = Switch_3_io_deqValid[2'h3:2'h3];
  assign T750 = {T751, io_deqValid_18};
  assign T751 = Switch_1_io_deqValid[1'h1:1'h1];
  assign T752 = {CU_1_io_deqValid, T753};
  assign T753 = {2'h0, CU_2_io_deqValid};
  assign T754 = {T761, T755};
  assign T755 = {T759, T756};
  assign T756 = {T758, T757};
  assign T757 = Switch_8_io_enqRdy[2'h2:2'h2];
  assign T758 = Switch_3_io_enqRdy[2'h3:2'h3];
  assign T759 = {T760, io_enqRdy_18};
  assign T760 = Switch_1_io_enqRdy[1'h1:1'h1];
  assign T761 = {CU_1_io_enqRdy, T762};
  assign T762 = {2'h3, CU_2_io_enqRdy};
  assign T763 = {CU_io_enqRdyOut, T764};
  assign T764 = {2'h3, CU_1_io_enqRdyOut};
  assign T765 = {T772, T766};
  assign T766 = {T770, T767};
  assign T767 = {T769, T768};
  assign T768 = Switch_7_io_deqValid[2'h2:2'h2];
  assign T769 = Switch_2_io_deqValid[2'h3:2'h3];
  assign T770 = {T771, io_deqValid_19};
  assign T771 = Switch_io_deqValid[1'h1:1'h1];
  assign T772 = {CU_io_deqValid, T773};
  assign T773 = {2'h0, CU_1_io_deqValid};
  assign T774 = {T781, T775};
  assign T775 = {T779, T776};
  assign T776 = {T778, T777};
  assign T777 = Switch_7_io_enqRdy[2'h2:2'h2];
  assign T778 = Switch_2_io_enqRdy[2'h3:2'h3];
  assign T779 = {T780, io_enqRdy_19};
  assign T780 = Switch_io_enqRdy[1'h1:1'h1];
  assign T781 = {CU_io_enqRdy, T782};
  assign T782 = {2'h3, CU_1_io_enqRdy};
  assign T783 = {3'h7, CU_io_enqRdyOut};
  assign T784 = {T789, T785};
  assign T785 = {1'h0, T786};
  assign T786 = {T788, T787};
  assign T787 = Switch_6_io_deqValid[2'h2:2'h2];
  assign T788 = Switch_1_io_deqValid[2'h3:2'h3];
  assign T789 = {3'h0, T790};
  assign T790 = {CU_io_deqValid, io_deqValid_0};
  assign T791 = {T796, T792};
  assign T792 = {1'h1, T793};
  assign T793 = {T795, T794};
  assign T794 = Switch_6_io_enqRdy[2'h2:2'h2];
  assign T795 = Switch_1_io_enqRdy[2'h3:2'h3];
  assign T796 = {3'h7, T797};
  assign T797 = {CU_io_enqRdy, io_enqRdy_0};
  assign T798 = {T802, T799};
  assign T799 = {T801, T800};
  assign T800 = Switch_35_io_deqValid[3'h6:3'h6];
  assign T801 = Switch_29_io_deqValid[3'h7:3'h7];
  assign T802 = {T804, T803};
  assign T803 = Switch_28_io_deqValid[3'h4:3'h4];
  assign T804 = Switch_34_io_deqValid[3'h5:3'h5];
  assign T805 = {T809, T806};
  assign T806 = {T808, T807};
  assign T807 = Switch_35_io_enqRdy[3'h6:3'h6];
  assign T808 = Switch_29_io_enqRdy[3'h7:3'h7];
  assign T809 = {T811, T810};
  assign T810 = Switch_28_io_enqRdy[3'h4:3'h4];
  assign T811 = Switch_34_io_enqRdy[3'h5:3'h5];
  assign T812 = {T816, T813};
  assign T813 = {T815, T814};
  assign T814 = Switch_34_io_deqValid[3'h6:3'h6];
  assign T815 = Switch_28_io_deqValid[3'h7:3'h7];
  assign T816 = {T818, T817};
  assign T817 = Switch_27_io_deqValid[3'h4:3'h4];
  assign T818 = Switch_33_io_deqValid[3'h5:3'h5];
  assign T819 = {T823, T820};
  assign T820 = {T822, T821};
  assign T821 = Switch_34_io_enqRdy[3'h6:3'h6];
  assign T822 = Switch_28_io_enqRdy[3'h7:3'h7];
  assign T823 = {T825, T824};
  assign T824 = Switch_27_io_enqRdy[3'h4:3'h4];
  assign T825 = Switch_33_io_enqRdy[3'h5:3'h5];
  assign T826 = {T830, T827};
  assign T827 = {T829, T828};
  assign T828 = Switch_33_io_deqValid[3'h6:3'h6];
  assign T829 = Switch_27_io_deqValid[3'h7:3'h7];
  assign T830 = {T832, T831};
  assign T831 = Switch_26_io_deqValid[3'h4:3'h4];
  assign T832 = Switch_32_io_deqValid[3'h5:3'h5];
  assign T833 = {T837, T834};
  assign T834 = {T836, T835};
  assign T835 = Switch_33_io_enqRdy[3'h6:3'h6];
  assign T836 = Switch_27_io_enqRdy[3'h7:3'h7];
  assign T837 = {T839, T838};
  assign T838 = Switch_26_io_enqRdy[3'h4:3'h4];
  assign T839 = Switch_32_io_enqRdy[3'h5:3'h5];
  assign T840 = {T844, T841};
  assign T841 = {T843, T842};
  assign T842 = Switch_32_io_deqValid[3'h6:3'h6];
  assign T843 = Switch_26_io_deqValid[3'h7:3'h7];
  assign T844 = {T846, T845};
  assign T845 = Switch_25_io_deqValid[3'h4:3'h4];
  assign T846 = Switch_31_io_deqValid[3'h5:3'h5];
  assign T847 = {T851, T848};
  assign T848 = {T850, T849};
  assign T849 = Switch_32_io_enqRdy[3'h6:3'h6];
  assign T850 = Switch_26_io_enqRdy[3'h7:3'h7];
  assign T851 = {T853, T852};
  assign T852 = Switch_25_io_enqRdy[3'h4:3'h4];
  assign T853 = Switch_31_io_enqRdy[3'h5:3'h5];
  assign T854 = {T858, T855};
  assign T855 = {T857, T856};
  assign T856 = Switch_31_io_deqValid[3'h6:3'h6];
  assign T857 = Switch_25_io_deqValid[3'h7:3'h7];
  assign T858 = {T860, T859};
  assign T859 = Switch_24_io_deqValid[3'h4:3'h4];
  assign T860 = Switch_30_io_deqValid[3'h5:3'h5];
  assign T861 = {T865, T862};
  assign T862 = {T864, T863};
  assign T863 = Switch_31_io_enqRdy[3'h6:3'h6];
  assign T864 = Switch_25_io_enqRdy[3'h7:3'h7];
  assign T865 = {T867, T866};
  assign T866 = Switch_24_io_enqRdy[3'h4:3'h4];
  assign T867 = Switch_30_io_enqRdy[3'h5:3'h5];
  assign T868 = {T872, T869};
  assign T869 = {T871, T870};
  assign T870 = Switch_29_io_deqValid[3'h6:3'h6];
  assign T871 = Switch_23_io_deqValid[3'h7:3'h7];
  assign T872 = {T874, T873};
  assign T873 = Switch_22_io_deqValid[3'h4:3'h4];
  assign T874 = Switch_28_io_deqValid[3'h5:3'h5];
  assign T875 = {T879, T876};
  assign T876 = {T878, T877};
  assign T877 = Switch_29_io_enqRdy[3'h6:3'h6];
  assign T878 = Switch_23_io_enqRdy[3'h7:3'h7];
  assign T879 = {T881, T880};
  assign T880 = Switch_22_io_enqRdy[3'h4:3'h4];
  assign T881 = Switch_28_io_enqRdy[3'h5:3'h5];
  assign T882 = {T886, T883};
  assign T883 = {T885, T884};
  assign T884 = Switch_28_io_deqValid[3'h6:3'h6];
  assign T885 = Switch_22_io_deqValid[3'h7:3'h7];
  assign T886 = {T888, T887};
  assign T887 = Switch_21_io_deqValid[3'h4:3'h4];
  assign T888 = Switch_27_io_deqValid[3'h5:3'h5];
  assign T889 = {T893, T890};
  assign T890 = {T892, T891};
  assign T891 = Switch_28_io_enqRdy[3'h6:3'h6];
  assign T892 = Switch_22_io_enqRdy[3'h7:3'h7];
  assign T893 = {T895, T894};
  assign T894 = Switch_21_io_enqRdy[3'h4:3'h4];
  assign T895 = Switch_27_io_enqRdy[3'h5:3'h5];
  assign T896 = {T900, T897};
  assign T897 = {T899, T898};
  assign T898 = Switch_27_io_deqValid[3'h6:3'h6];
  assign T899 = Switch_21_io_deqValid[3'h7:3'h7];
  assign T900 = {T902, T901};
  assign T901 = Switch_20_io_deqValid[3'h4:3'h4];
  assign T902 = Switch_26_io_deqValid[3'h5:3'h5];
  assign T903 = {T907, T904};
  assign T904 = {T906, T905};
  assign T905 = Switch_27_io_enqRdy[3'h6:3'h6];
  assign T906 = Switch_21_io_enqRdy[3'h7:3'h7];
  assign T907 = {T909, T908};
  assign T908 = Switch_20_io_enqRdy[3'h4:3'h4];
  assign T909 = Switch_26_io_enqRdy[3'h5:3'h5];
  assign T910 = {T914, T911};
  assign T911 = {T913, T912};
  assign T912 = Switch_26_io_deqValid[3'h6:3'h6];
  assign T913 = Switch_20_io_deqValid[3'h7:3'h7];
  assign T914 = {T916, T915};
  assign T915 = Switch_19_io_deqValid[3'h4:3'h4];
  assign T916 = Switch_25_io_deqValid[3'h5:3'h5];
  assign T917 = {T921, T918};
  assign T918 = {T920, T919};
  assign T919 = Switch_26_io_enqRdy[3'h6:3'h6];
  assign T920 = Switch_20_io_enqRdy[3'h7:3'h7];
  assign T921 = {T923, T922};
  assign T922 = Switch_19_io_enqRdy[3'h4:3'h4];
  assign T923 = Switch_25_io_enqRdy[3'h5:3'h5];
  assign T924 = {T928, T925};
  assign T925 = {T927, T926};
  assign T926 = Switch_25_io_deqValid[3'h6:3'h6];
  assign T927 = Switch_19_io_deqValid[3'h7:3'h7];
  assign T928 = {T930, T929};
  assign T929 = Switch_18_io_deqValid[3'h4:3'h4];
  assign T930 = Switch_24_io_deqValid[3'h5:3'h5];
  assign T931 = {T935, T932};
  assign T932 = {T934, T933};
  assign T933 = Switch_25_io_enqRdy[3'h6:3'h6];
  assign T934 = Switch_19_io_enqRdy[3'h7:3'h7];
  assign T935 = {T937, T936};
  assign T936 = Switch_18_io_enqRdy[3'h4:3'h4];
  assign T937 = Switch_24_io_enqRdy[3'h5:3'h5];
  assign T938 = {T942, T939};
  assign T939 = {T941, T940};
  assign T940 = Switch_23_io_deqValid[3'h6:3'h6];
  assign T941 = Switch_17_io_deqValid[3'h7:3'h7];
  assign T942 = {T944, T943};
  assign T943 = Switch_16_io_deqValid[3'h4:3'h4];
  assign T944 = Switch_22_io_deqValid[3'h5:3'h5];
  assign T945 = {T949, T946};
  assign T946 = {T948, T947};
  assign T947 = Switch_23_io_enqRdy[3'h6:3'h6];
  assign T948 = Switch_17_io_enqRdy[3'h7:3'h7];
  assign T949 = {T951, T950};
  assign T950 = Switch_16_io_enqRdy[3'h4:3'h4];
  assign T951 = Switch_22_io_enqRdy[3'h5:3'h5];
  assign T952 = {T956, T953};
  assign T953 = {T955, T954};
  assign T954 = Switch_22_io_deqValid[3'h6:3'h6];
  assign T955 = Switch_16_io_deqValid[3'h7:3'h7];
  assign T956 = {T958, T957};
  assign T957 = Switch_15_io_deqValid[3'h4:3'h4];
  assign T958 = Switch_21_io_deqValid[3'h5:3'h5];
  assign T959 = {T963, T960};
  assign T960 = {T962, T961};
  assign T961 = Switch_22_io_enqRdy[3'h6:3'h6];
  assign T962 = Switch_16_io_enqRdy[3'h7:3'h7];
  assign T963 = {T965, T964};
  assign T964 = Switch_15_io_enqRdy[3'h4:3'h4];
  assign T965 = Switch_21_io_enqRdy[3'h5:3'h5];
  assign T966 = {T970, T967};
  assign T967 = {T969, T968};
  assign T968 = Switch_21_io_deqValid[3'h6:3'h6];
  assign T969 = Switch_15_io_deqValid[3'h7:3'h7];
  assign T970 = {T972, T971};
  assign T971 = Switch_14_io_deqValid[3'h4:3'h4];
  assign T972 = Switch_20_io_deqValid[3'h5:3'h5];
  assign T973 = {T977, T974};
  assign T974 = {T976, T975};
  assign T975 = Switch_21_io_enqRdy[3'h6:3'h6];
  assign T976 = Switch_15_io_enqRdy[3'h7:3'h7];
  assign T977 = {T979, T978};
  assign T978 = Switch_14_io_enqRdy[3'h4:3'h4];
  assign T979 = Switch_20_io_enqRdy[3'h5:3'h5];
  assign T980 = {T984, T981};
  assign T981 = {T983, T982};
  assign T982 = Switch_20_io_deqValid[3'h6:3'h6];
  assign T983 = Switch_14_io_deqValid[3'h7:3'h7];
  assign T984 = {T986, T985};
  assign T985 = Switch_13_io_deqValid[3'h4:3'h4];
  assign T986 = Switch_19_io_deqValid[3'h5:3'h5];
  assign T987 = {T991, T988};
  assign T988 = {T990, T989};
  assign T989 = Switch_20_io_enqRdy[3'h6:3'h6];
  assign T990 = Switch_14_io_enqRdy[3'h7:3'h7];
  assign T991 = {T993, T992};
  assign T992 = Switch_13_io_enqRdy[3'h4:3'h4];
  assign T993 = Switch_19_io_enqRdy[3'h5:3'h5];
  assign T994 = {T998, T995};
  assign T995 = {T997, T996};
  assign T996 = Switch_19_io_deqValid[3'h6:3'h6];
  assign T997 = Switch_13_io_deqValid[3'h7:3'h7];
  assign T998 = {T1000, T999};
  assign T999 = Switch_12_io_deqValid[3'h4:3'h4];
  assign T1000 = Switch_18_io_deqValid[3'h5:3'h5];
  assign T1001 = {T1005, T1002};
  assign T1002 = {T1004, T1003};
  assign T1003 = Switch_19_io_enqRdy[3'h6:3'h6];
  assign T1004 = Switch_13_io_enqRdy[3'h7:3'h7];
  assign T1005 = {T1007, T1006};
  assign T1006 = Switch_12_io_enqRdy[3'h4:3'h4];
  assign T1007 = Switch_18_io_enqRdy[3'h5:3'h5];
  assign T1008 = {T1012, T1009};
  assign T1009 = {T1011, T1010};
  assign T1010 = Switch_17_io_deqValid[3'h6:3'h6];
  assign T1011 = Switch_11_io_deqValid[3'h7:3'h7];
  assign T1012 = {T1014, T1013};
  assign T1013 = Switch_10_io_deqValid[3'h4:3'h4];
  assign T1014 = Switch_16_io_deqValid[3'h5:3'h5];
  assign T1015 = {T1019, T1016};
  assign T1016 = {T1018, T1017};
  assign T1017 = Switch_17_io_enqRdy[3'h6:3'h6];
  assign T1018 = Switch_11_io_enqRdy[3'h7:3'h7];
  assign T1019 = {T1021, T1020};
  assign T1020 = Switch_10_io_enqRdy[3'h4:3'h4];
  assign T1021 = Switch_16_io_enqRdy[3'h5:3'h5];
  assign T1022 = {T1026, T1023};
  assign T1023 = {T1025, T1024};
  assign T1024 = Switch_16_io_deqValid[3'h6:3'h6];
  assign T1025 = Switch_10_io_deqValid[3'h7:3'h7];
  assign T1026 = {T1028, T1027};
  assign T1027 = Switch_9_io_deqValid[3'h4:3'h4];
  assign T1028 = Switch_15_io_deqValid[3'h5:3'h5];
  assign T1029 = {T1033, T1030};
  assign T1030 = {T1032, T1031};
  assign T1031 = Switch_16_io_enqRdy[3'h6:3'h6];
  assign T1032 = Switch_10_io_enqRdy[3'h7:3'h7];
  assign T1033 = {T1035, T1034};
  assign T1034 = Switch_9_io_enqRdy[3'h4:3'h4];
  assign T1035 = Switch_15_io_enqRdy[3'h5:3'h5];
  assign T1036 = {T1040, T1037};
  assign T1037 = {T1039, T1038};
  assign T1038 = Switch_15_io_deqValid[3'h6:3'h6];
  assign T1039 = Switch_9_io_deqValid[3'h7:3'h7];
  assign T1040 = {T1042, T1041};
  assign T1041 = Switch_8_io_deqValid[3'h4:3'h4];
  assign T1042 = Switch_14_io_deqValid[3'h5:3'h5];
  assign T1043 = {T1047, T1044};
  assign T1044 = {T1046, T1045};
  assign T1045 = Switch_15_io_enqRdy[3'h6:3'h6];
  assign T1046 = Switch_9_io_enqRdy[3'h7:3'h7];
  assign T1047 = {T1049, T1048};
  assign T1048 = Switch_8_io_enqRdy[3'h4:3'h4];
  assign T1049 = Switch_14_io_enqRdy[3'h5:3'h5];
  assign T1050 = {T1054, T1051};
  assign T1051 = {T1053, T1052};
  assign T1052 = Switch_14_io_deqValid[3'h6:3'h6];
  assign T1053 = Switch_8_io_deqValid[3'h7:3'h7];
  assign T1054 = {T1056, T1055};
  assign T1055 = Switch_7_io_deqValid[3'h4:3'h4];
  assign T1056 = Switch_13_io_deqValid[3'h5:3'h5];
  assign T1057 = {T1061, T1058};
  assign T1058 = {T1060, T1059};
  assign T1059 = Switch_14_io_enqRdy[3'h6:3'h6];
  assign T1060 = Switch_8_io_enqRdy[3'h7:3'h7];
  assign T1061 = {T1063, T1062};
  assign T1062 = Switch_7_io_enqRdy[3'h4:3'h4];
  assign T1063 = Switch_13_io_enqRdy[3'h5:3'h5];
  assign T1064 = {T1068, T1065};
  assign T1065 = {T1067, T1066};
  assign T1066 = Switch_13_io_deqValid[3'h6:3'h6];
  assign T1067 = Switch_7_io_deqValid[3'h7:3'h7];
  assign T1068 = {T1070, T1069};
  assign T1069 = Switch_6_io_deqValid[3'h4:3'h4];
  assign T1070 = Switch_12_io_deqValid[3'h5:3'h5];
  assign T1071 = {T1075, T1072};
  assign T1072 = {T1074, T1073};
  assign T1073 = Switch_13_io_enqRdy[3'h6:3'h6];
  assign T1074 = Switch_7_io_enqRdy[3'h7:3'h7];
  assign T1075 = {T1077, T1076};
  assign T1076 = Switch_6_io_enqRdy[3'h4:3'h4];
  assign T1077 = Switch_12_io_enqRdy[3'h5:3'h5];
  assign T1078 = {T1082, T1079};
  assign T1079 = {T1081, T1080};
  assign T1080 = Switch_11_io_deqValid[3'h6:3'h6];
  assign T1081 = Switch_5_io_deqValid[3'h7:3'h7];
  assign T1082 = {T1084, T1083};
  assign T1083 = Switch_4_io_deqValid[3'h4:3'h4];
  assign T1084 = Switch_10_io_deqValid[3'h5:3'h5];
  assign T1085 = {T1089, T1086};
  assign T1086 = {T1088, T1087};
  assign T1087 = Switch_11_io_enqRdy[3'h6:3'h6];
  assign T1088 = Switch_5_io_enqRdy[3'h7:3'h7];
  assign T1089 = {T1091, T1090};
  assign T1090 = Switch_4_io_enqRdy[3'h4:3'h4];
  assign T1091 = Switch_10_io_enqRdy[3'h5:3'h5];
  assign T1092 = {T1096, T1093};
  assign T1093 = {T1095, T1094};
  assign T1094 = Switch_10_io_deqValid[3'h6:3'h6];
  assign T1095 = Switch_4_io_deqValid[3'h7:3'h7];
  assign T1096 = {T1098, T1097};
  assign T1097 = Switch_3_io_deqValid[3'h4:3'h4];
  assign T1098 = Switch_9_io_deqValid[3'h5:3'h5];
  assign T1099 = {T1103, T1100};
  assign T1100 = {T1102, T1101};
  assign T1101 = Switch_10_io_enqRdy[3'h6:3'h6];
  assign T1102 = Switch_4_io_enqRdy[3'h7:3'h7];
  assign T1103 = {T1105, T1104};
  assign T1104 = Switch_3_io_enqRdy[3'h4:3'h4];
  assign T1105 = Switch_9_io_enqRdy[3'h5:3'h5];
  assign T1106 = {T1110, T1107};
  assign T1107 = {T1109, T1108};
  assign T1108 = Switch_9_io_deqValid[3'h6:3'h6];
  assign T1109 = Switch_3_io_deqValid[3'h7:3'h7];
  assign T1110 = {T1112, T1111};
  assign T1111 = Switch_2_io_deqValid[3'h4:3'h4];
  assign T1112 = Switch_8_io_deqValid[3'h5:3'h5];
  assign T1113 = {T1117, T1114};
  assign T1114 = {T1116, T1115};
  assign T1115 = Switch_9_io_enqRdy[3'h6:3'h6];
  assign T1116 = Switch_3_io_enqRdy[3'h7:3'h7];
  assign T1117 = {T1119, T1118};
  assign T1118 = Switch_2_io_enqRdy[3'h4:3'h4];
  assign T1119 = Switch_8_io_enqRdy[3'h5:3'h5];
  assign T1120 = {T1124, T1121};
  assign T1121 = {T1123, T1122};
  assign T1122 = Switch_8_io_deqValid[3'h6:3'h6];
  assign T1123 = Switch_2_io_deqValid[3'h7:3'h7];
  assign T1124 = {T1126, T1125};
  assign T1125 = Switch_1_io_deqValid[3'h4:3'h4];
  assign T1126 = Switch_7_io_deqValid[3'h5:3'h5];
  assign T1127 = {T1131, T1128};
  assign T1128 = {T1130, T1129};
  assign T1129 = Switch_8_io_enqRdy[3'h6:3'h6];
  assign T1130 = Switch_2_io_enqRdy[3'h7:3'h7];
  assign T1131 = {T1133, T1132};
  assign T1132 = Switch_1_io_enqRdy[3'h4:3'h4];
  assign T1133 = Switch_7_io_enqRdy[3'h5:3'h5];
  assign T1134 = {T1138, T1135};
  assign T1135 = {T1137, T1136};
  assign T1136 = Switch_7_io_deqValid[3'h6:3'h6];
  assign T1137 = Switch_1_io_deqValid[3'h7:3'h7];
  assign T1138 = {T1140, T1139};
  assign T1139 = Switch_io_deqValid[3'h4:3'h4];
  assign T1140 = Switch_6_io_deqValid[3'h5:3'h5];
  assign T1141 = {T1145, T1142};
  assign T1142 = {T1144, T1143};
  assign T1143 = Switch_7_io_enqRdy[3'h6:3'h6];
  assign T1144 = Switch_1_io_enqRdy[3'h7:3'h7];
  assign T1145 = {T1147, T1146};
  assign T1146 = Switch_io_enqRdy[3'h4:3'h4];
  assign T1147 = Switch_6_io_enqRdy[3'h5:3'h5];
  assign io_enqValid_0 = T1148;
  assign T1148 = Switch_io_deqValid[2'h3:2'h3];
  assign io_enqValid_1 = T1149;
  assign T1149 = Switch_6_io_deqValid[2'h3:2'h3];
  assign io_enqValid_2 = T1150;
  assign T1150 = Switch_12_io_deqValid[2'h3:2'h3];
  assign io_enqValid_3 = T1151;
  assign T1151 = Switch_18_io_deqValid[2'h3:2'h3];
  assign io_enqValid_4 = T1152;
  assign T1152 = Switch_24_io_deqValid[2'h3:2'h3];
  assign io_enqValid_5 = T1153;
  assign T1153 = Switch_30_io_deqValid[2'h3:2'h3];
  assign io_enqValid_6 = T1154;
  assign T1154 = Switch_31_io_deqValid[1'h0:1'h0];
  assign io_enqValid_7 = T1155;
  assign T1155 = Switch_32_io_deqValid[1'h0:1'h0];
  assign io_enqValid_8 = T1156;
  assign T1156 = Switch_33_io_deqValid[1'h0:1'h0];
  assign io_enqValid_9 = T1157;
  assign T1157 = Switch_34_io_deqValid[1'h0:1'h0];
  assign io_enqValid_10 = T1158;
  assign T1158 = Switch_35_io_deqValid[1'h1:1'h1];
  assign io_enqValid_11 = T1159;
  assign T1159 = Switch_29_io_deqValid[1'h1:1'h1];
  assign io_enqValid_12 = T1160;
  assign T1160 = Switch_23_io_deqValid[1'h1:1'h1];
  assign io_enqValid_13 = T1161;
  assign T1161 = Switch_17_io_deqValid[1'h1:1'h1];
  assign io_enqValid_14 = T1162;
  assign T1162 = Switch_11_io_deqValid[1'h1:1'h1];
  assign io_enqValid_15 = T1163;
  assign T1163 = Switch_5_io_deqValid[1'h1:1'h1];
  assign io_enqValid_16 = T1164;
  assign T1164 = Switch_4_io_deqValid[2'h2:2'h2];
  assign io_enqValid_17 = T1165;
  assign T1165 = Switch_3_io_deqValid[2'h2:2'h2];
  assign io_enqValid_18 = T1166;
  assign T1166 = Switch_2_io_deqValid[2'h2:2'h2];
  assign io_enqValid_19 = T1167;
  assign T1167 = Switch_1_io_deqValid[2'h2:2'h2];
  assign io_deqRdy_0 = T1168;
  assign T1168 = Switch_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_1 = T1169;
  assign T1169 = Switch_6_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_2 = T1170;
  assign T1170 = Switch_12_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_3 = T1171;
  assign T1171 = Switch_18_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_4 = T1172;
  assign T1172 = Switch_24_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_5 = T1173;
  assign T1173 = Switch_30_io_enqRdy[2'h3:2'h3];
  assign io_deqRdy_6 = T1174;
  assign T1174 = Switch_31_io_enqRdy[1'h0:1'h0];
  assign io_deqRdy_7 = T1175;
  assign T1175 = Switch_32_io_enqRdy[1'h0:1'h0];
  assign io_deqRdy_8 = T1176;
  assign T1176 = Switch_33_io_enqRdy[1'h0:1'h0];
  assign io_deqRdy_9 = T1177;
  assign T1177 = Switch_34_io_enqRdy[1'h0:1'h0];
  assign io_deqRdy_10 = T1178;
  assign T1178 = Switch_35_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_11 = T1179;
  assign T1179 = Switch_29_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_12 = T1180;
  assign T1180 = Switch_23_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_13 = T1181;
  assign T1181 = Switch_17_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_14 = T1182;
  assign T1182 = Switch_11_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_15 = T1183;
  assign T1183 = Switch_5_io_enqRdy[1'h1:1'h1];
  assign io_deqRdy_16 = T1184;
  assign T1184 = Switch_4_io_enqRdy[2'h2:2'h2];
  assign io_deqRdy_17 = T1185;
  assign T1185 = Switch_3_io_enqRdy[2'h2:2'h2];
  assign io_deqRdy_18 = T1186;
  assign T1186 = Switch_2_io_enqRdy[2'h2:2'h2];
  assign io_deqRdy_19 = T1187;
  assign T1187 = Switch_1_io_enqRdy[2'h2:2'h2];
  assign io_outData_0 = Switch_io_outPort_3;
  assign io_outData_1 = Switch_6_io_outPort_3;
  assign io_outData_2 = Switch_12_io_outPort_3;
  assign io_outData_3 = Switch_18_io_outPort_3;
  assign io_outData_4 = Switch_24_io_outPort_3;
  assign io_outData_5 = Switch_30_io_outPort_3;
  assign io_outData_6 = Switch_31_io_outPort_0;
  assign io_outData_7 = Switch_32_io_outPort_0;
  assign io_outData_8 = Switch_33_io_outPort_0;
  assign io_outData_9 = Switch_34_io_outPort_0;
  assign io_outData_10 = Switch_35_io_outPort_1;
  assign io_outData_11 = Switch_29_io_outPort_1;
  assign io_outData_12 = Switch_23_io_outPort_1;
  assign io_outData_13 = Switch_17_io_outPort_1;
  assign io_outData_14 = Switch_11_io_outPort_1;
  assign io_outData_15 = Switch_5_io_outPort_1;
  assign io_outData_16 = Switch_4_io_outPort_2;
  assign io_outData_17 = Switch_3_io_outPort_2;
  assign io_outData_18 = Switch_2_io_outPort_2;
  assign io_outData_19 = Switch_1_io_outPort_2;
  CU CU(.clk(clk), .reset(reset),
       .io_in_3( Switch_6_io_outPort_5 ),
       .io_in_2( Switch_io_outPort_4 ),
       .io_in_1( Switch_1_io_outPort_7 ),
       .io_in_0( Switch_7_io_outPort_6 ),
       .io_out( CU_io_out ),
       .io_inConfig( Switch_io_outCUConfig ),
       .io_enqRdy( CU_io_enqRdy ),
       .io_deqRdy( T1141 ),
       .io_enqValid( T1134 ),
       .io_deqValid( CU_io_deqValid ),
       .io_enqRdyOut( CU_io_enqRdyOut )
  );
  CU CU_1(.clk(clk), .reset(reset),
       .io_in_3( Switch_7_io_outPort_5 ),
       .io_in_2( Switch_1_io_outPort_4 ),
       .io_in_1( Switch_2_io_outPort_7 ),
       .io_in_0( Switch_8_io_outPort_6 ),
       .io_out( CU_1_io_out ),
       .io_inConfig( Switch_1_io_outCUConfig ),
       .io_enqRdy( CU_1_io_enqRdy ),
       .io_deqRdy( T1127 ),
       .io_enqValid( T1120 ),
       .io_deqValid( CU_1_io_deqValid ),
       .io_enqRdyOut( CU_1_io_enqRdyOut )
  );
  CU CU_2(.clk(clk), .reset(reset),
       .io_in_3( Switch_8_io_outPort_5 ),
       .io_in_2( Switch_2_io_outPort_4 ),
       .io_in_1( Switch_3_io_outPort_7 ),
       .io_in_0( Switch_9_io_outPort_6 ),
       .io_out( CU_2_io_out ),
       .io_inConfig( Switch_2_io_outCUConfig ),
       .io_enqRdy( CU_2_io_enqRdy ),
       .io_deqRdy( T1113 ),
       .io_enqValid( T1106 ),
       .io_deqValid( CU_2_io_deqValid ),
       .io_enqRdyOut( CU_2_io_enqRdyOut )
  );
  CU CU_3(.clk(clk), .reset(reset),
       .io_in_3( Switch_9_io_outPort_5 ),
       .io_in_2( Switch_3_io_outPort_4 ),
       .io_in_1( Switch_4_io_outPort_7 ),
       .io_in_0( Switch_10_io_outPort_6 ),
       .io_out( CU_3_io_out ),
       .io_inConfig( Switch_3_io_outCUConfig ),
       .io_enqRdy( CU_3_io_enqRdy ),
       .io_deqRdy( T1099 ),
       .io_enqValid( T1092 ),
       .io_deqValid( CU_3_io_deqValid ),
       .io_enqRdyOut( CU_3_io_enqRdyOut )
  );
  CU CU_4(.clk(clk), .reset(reset),
       .io_in_3( Switch_10_io_outPort_5 ),
       .io_in_2( Switch_4_io_outPort_4 ),
       .io_in_1( Switch_5_io_outPort_7 ),
       .io_in_0( Switch_11_io_outPort_6 ),
       .io_out( CU_4_io_out ),
       .io_inConfig( Switch_4_io_outCUConfig ),
       .io_enqRdy( CU_4_io_enqRdy ),
       .io_deqRdy( T1085 ),
       .io_enqValid( T1078 ),
       .io_deqValid( CU_4_io_deqValid ),
       .io_enqRdyOut( CU_4_io_enqRdyOut )
  );
  CU CU_5(.clk(clk), .reset(reset),
       .io_in_3( Switch_12_io_outPort_5 ),
       .io_in_2( Switch_6_io_outPort_4 ),
       .io_in_1( Switch_7_io_outPort_7 ),
       .io_in_0( Switch_13_io_outPort_6 ),
       .io_out( CU_5_io_out ),
       .io_inConfig( Switch_6_io_outCUConfig ),
       .io_enqRdy( CU_5_io_enqRdy ),
       .io_deqRdy( T1071 ),
       .io_enqValid( T1064 ),
       .io_deqValid( CU_5_io_deqValid ),
       .io_enqRdyOut( CU_5_io_enqRdyOut )
  );
  CU CU_6(.clk(clk), .reset(reset),
       .io_in_3( Switch_13_io_outPort_5 ),
       .io_in_2( Switch_7_io_outPort_4 ),
       .io_in_1( Switch_8_io_outPort_7 ),
       .io_in_0( Switch_14_io_outPort_6 ),
       .io_out( CU_6_io_out ),
       .io_inConfig( Switch_7_io_outCUConfig ),
       .io_enqRdy( CU_6_io_enqRdy ),
       .io_deqRdy( T1057 ),
       .io_enqValid( T1050 ),
       .io_deqValid( CU_6_io_deqValid ),
       .io_enqRdyOut( CU_6_io_enqRdyOut )
  );
  CU CU_7(.clk(clk), .reset(reset),
       .io_in_3( Switch_14_io_outPort_5 ),
       .io_in_2( Switch_8_io_outPort_4 ),
       .io_in_1( Switch_9_io_outPort_7 ),
       .io_in_0( Switch_15_io_outPort_6 ),
       .io_out( CU_7_io_out ),
       .io_inConfig( Switch_8_io_outCUConfig ),
       .io_enqRdy( CU_7_io_enqRdy ),
       .io_deqRdy( T1043 ),
       .io_enqValid( T1036 ),
       .io_deqValid( CU_7_io_deqValid ),
       .io_enqRdyOut( CU_7_io_enqRdyOut )
  );
  CU CU_8(.clk(clk), .reset(reset),
       .io_in_3( Switch_15_io_outPort_5 ),
       .io_in_2( Switch_9_io_outPort_4 ),
       .io_in_1( Switch_10_io_outPort_7 ),
       .io_in_0( Switch_16_io_outPort_6 ),
       .io_out( CU_8_io_out ),
       .io_inConfig( Switch_9_io_outCUConfig ),
       .io_enqRdy( CU_8_io_enqRdy ),
       .io_deqRdy( T1029 ),
       .io_enqValid( T1022 ),
       .io_deqValid( CU_8_io_deqValid ),
       .io_enqRdyOut( CU_8_io_enqRdyOut )
  );
  CU CU_9(.clk(clk), .reset(reset),
       .io_in_3( Switch_16_io_outPort_5 ),
       .io_in_2( Switch_10_io_outPort_4 ),
       .io_in_1( Switch_11_io_outPort_7 ),
       .io_in_0( Switch_17_io_outPort_6 ),
       .io_out( CU_9_io_out ),
       .io_inConfig( Switch_10_io_outCUConfig ),
       .io_enqRdy( CU_9_io_enqRdy ),
       .io_deqRdy( T1015 ),
       .io_enqValid( T1008 ),
       .io_deqValid( CU_9_io_deqValid ),
       .io_enqRdyOut( CU_9_io_enqRdyOut )
  );
  CU CU_10(.clk(clk), .reset(reset),
       .io_in_3( Switch_18_io_outPort_5 ),
       .io_in_2( Switch_12_io_outPort_4 ),
       .io_in_1( Switch_13_io_outPort_7 ),
       .io_in_0( Switch_19_io_outPort_6 ),
       .io_out( CU_10_io_out ),
       .io_inConfig( Switch_12_io_outCUConfig ),
       .io_enqRdy( CU_10_io_enqRdy ),
       .io_deqRdy( T1001 ),
       .io_enqValid( T994 ),
       .io_deqValid( CU_10_io_deqValid ),
       .io_enqRdyOut( CU_10_io_enqRdyOut )
  );
  CU CU_11(.clk(clk), .reset(reset),
       .io_in_3( Switch_19_io_outPort_5 ),
       .io_in_2( Switch_13_io_outPort_4 ),
       .io_in_1( Switch_14_io_outPort_7 ),
       .io_in_0( Switch_20_io_outPort_6 ),
       .io_out( CU_11_io_out ),
       .io_inConfig( Switch_13_io_outCUConfig ),
       .io_enqRdy( CU_11_io_enqRdy ),
       .io_deqRdy( T987 ),
       .io_enqValid( T980 ),
       .io_deqValid( CU_11_io_deqValid ),
       .io_enqRdyOut( CU_11_io_enqRdyOut )
  );
  CU CU_12(.clk(clk), .reset(reset),
       .io_in_3( Switch_20_io_outPort_5 ),
       .io_in_2( Switch_14_io_outPort_4 ),
       .io_in_1( Switch_15_io_outPort_7 ),
       .io_in_0( Switch_21_io_outPort_6 ),
       .io_out( CU_12_io_out ),
       .io_inConfig( Switch_14_io_outCUConfig ),
       .io_enqRdy( CU_12_io_enqRdy ),
       .io_deqRdy( T973 ),
       .io_enqValid( T966 ),
       .io_deqValid( CU_12_io_deqValid ),
       .io_enqRdyOut( CU_12_io_enqRdyOut )
  );
  CU CU_13(.clk(clk), .reset(reset),
       .io_in_3( Switch_21_io_outPort_5 ),
       .io_in_2( Switch_15_io_outPort_4 ),
       .io_in_1( Switch_16_io_outPort_7 ),
       .io_in_0( Switch_22_io_outPort_6 ),
       .io_out( CU_13_io_out ),
       .io_inConfig( Switch_15_io_outCUConfig ),
       .io_enqRdy( CU_13_io_enqRdy ),
       .io_deqRdy( T959 ),
       .io_enqValid( T952 ),
       .io_deqValid( CU_13_io_deqValid ),
       .io_enqRdyOut( CU_13_io_enqRdyOut )
  );
  CU CU_14(.clk(clk), .reset(reset),
       .io_in_3( Switch_22_io_outPort_5 ),
       .io_in_2( Switch_16_io_outPort_4 ),
       .io_in_1( Switch_17_io_outPort_7 ),
       .io_in_0( Switch_23_io_outPort_6 ),
       .io_out( CU_14_io_out ),
       .io_inConfig( Switch_16_io_outCUConfig ),
       .io_enqRdy( CU_14_io_enqRdy ),
       .io_deqRdy( T945 ),
       .io_enqValid( T938 ),
       .io_deqValid( CU_14_io_deqValid ),
       .io_enqRdyOut( CU_14_io_enqRdyOut )
  );
  CU CU_15(.clk(clk), .reset(reset),
       .io_in_3( Switch_24_io_outPort_5 ),
       .io_in_2( Switch_18_io_outPort_4 ),
       .io_in_1( Switch_19_io_outPort_7 ),
       .io_in_0( Switch_25_io_outPort_6 ),
       .io_out( CU_15_io_out ),
       .io_inConfig( Switch_18_io_outCUConfig ),
       .io_enqRdy( CU_15_io_enqRdy ),
       .io_deqRdy( T931 ),
       .io_enqValid( T924 ),
       .io_deqValid( CU_15_io_deqValid ),
       .io_enqRdyOut( CU_15_io_enqRdyOut )
  );
  CU CU_16(.clk(clk), .reset(reset),
       .io_in_3( Switch_25_io_outPort_5 ),
       .io_in_2( Switch_19_io_outPort_4 ),
       .io_in_1( Switch_20_io_outPort_7 ),
       .io_in_0( Switch_26_io_outPort_6 ),
       .io_out( CU_16_io_out ),
       .io_inConfig( Switch_19_io_outCUConfig ),
       .io_enqRdy( CU_16_io_enqRdy ),
       .io_deqRdy( T917 ),
       .io_enqValid( T910 ),
       .io_deqValid( CU_16_io_deqValid ),
       .io_enqRdyOut( CU_16_io_enqRdyOut )
  );
  CU CU_17(.clk(clk), .reset(reset),
       .io_in_3( Switch_26_io_outPort_5 ),
       .io_in_2( Switch_20_io_outPort_4 ),
       .io_in_1( Switch_21_io_outPort_7 ),
       .io_in_0( Switch_27_io_outPort_6 ),
       .io_out( CU_17_io_out ),
       .io_inConfig( Switch_20_io_outCUConfig ),
       .io_enqRdy( CU_17_io_enqRdy ),
       .io_deqRdy( T903 ),
       .io_enqValid( T896 ),
       .io_deqValid( CU_17_io_deqValid ),
       .io_enqRdyOut( CU_17_io_enqRdyOut )
  );
  CU CU_18(.clk(clk), .reset(reset),
       .io_in_3( Switch_27_io_outPort_5 ),
       .io_in_2( Switch_21_io_outPort_4 ),
       .io_in_1( Switch_22_io_outPort_7 ),
       .io_in_0( Switch_28_io_outPort_6 ),
       .io_out( CU_18_io_out ),
       .io_inConfig( Switch_21_io_outCUConfig ),
       .io_enqRdy( CU_18_io_enqRdy ),
       .io_deqRdy( T889 ),
       .io_enqValid( T882 ),
       .io_deqValid( CU_18_io_deqValid ),
       .io_enqRdyOut( CU_18_io_enqRdyOut )
  );
  CU CU_19(.clk(clk), .reset(reset),
       .io_in_3( Switch_28_io_outPort_5 ),
       .io_in_2( Switch_22_io_outPort_4 ),
       .io_in_1( Switch_23_io_outPort_7 ),
       .io_in_0( Switch_29_io_outPort_6 ),
       .io_out( CU_19_io_out ),
       .io_inConfig( Switch_22_io_outCUConfig ),
       .io_enqRdy( CU_19_io_enqRdy ),
       .io_deqRdy( T875 ),
       .io_enqValid( T868 ),
       .io_deqValid( CU_19_io_deqValid ),
       .io_enqRdyOut( CU_19_io_enqRdyOut )
  );
  CU CU_20(.clk(clk), .reset(reset),
       .io_in_3( Switch_30_io_outPort_5 ),
       .io_in_2( Switch_24_io_outPort_4 ),
       .io_in_1( Switch_25_io_outPort_7 ),
       .io_in_0( Switch_31_io_outPort_6 ),
       .io_out( CU_20_io_out ),
       .io_inConfig( Switch_24_io_outCUConfig ),
       .io_enqRdy( CU_20_io_enqRdy ),
       .io_deqRdy( T861 ),
       .io_enqValid( T854 ),
       .io_deqValid( CU_20_io_deqValid ),
       .io_enqRdyOut( CU_20_io_enqRdyOut )
  );
  CU CU_21(.clk(clk), .reset(reset),
       .io_in_3( Switch_31_io_outPort_5 ),
       .io_in_2( Switch_25_io_outPort_4 ),
       .io_in_1( Switch_26_io_outPort_7 ),
       .io_in_0( Switch_32_io_outPort_6 ),
       .io_out( CU_21_io_out ),
       .io_inConfig( Switch_25_io_outCUConfig ),
       .io_enqRdy( CU_21_io_enqRdy ),
       .io_deqRdy( T847 ),
       .io_enqValid( T840 ),
       .io_deqValid( CU_21_io_deqValid ),
       .io_enqRdyOut( CU_21_io_enqRdyOut )
  );
  CU CU_22(.clk(clk), .reset(reset),
       .io_in_3( Switch_32_io_outPort_5 ),
       .io_in_2( Switch_26_io_outPort_4 ),
       .io_in_1( Switch_27_io_outPort_7 ),
       .io_in_0( Switch_33_io_outPort_6 ),
       .io_out( CU_22_io_out ),
       .io_inConfig( Switch_26_io_outCUConfig ),
       .io_enqRdy( CU_22_io_enqRdy ),
       .io_deqRdy( T833 ),
       .io_enqValid( T826 ),
       .io_deqValid( CU_22_io_deqValid ),
       .io_enqRdyOut( CU_22_io_enqRdyOut )
  );
  CU CU_23(.clk(clk), .reset(reset),
       .io_in_3( Switch_33_io_outPort_5 ),
       .io_in_2( Switch_27_io_outPort_4 ),
       .io_in_1( Switch_28_io_outPort_7 ),
       .io_in_0( Switch_34_io_outPort_6 ),
       .io_out( CU_23_io_out ),
       .io_inConfig( Switch_27_io_outCUConfig ),
       .io_enqRdy( CU_23_io_enqRdy ),
       .io_deqRdy( T819 ),
       .io_enqValid( T812 ),
       .io_deqValid( CU_23_io_deqValid ),
       .io_enqRdyOut( CU_23_io_enqRdyOut )
  );
  CU CU_24(.clk(clk), .reset(reset),
       .io_in_3( Switch_34_io_outPort_5 ),
       .io_in_2( Switch_28_io_outPort_4 ),
       .io_in_1( Switch_29_io_outPort_7 ),
       .io_in_0( Switch_35_io_outPort_6 ),
       .io_out( CU_24_io_out ),
       .io_inConfig( Switch_28_io_outCUConfig ),
       .io_enqRdy( CU_24_io_enqRdy ),
       .io_deqRdy( T805 ),
       .io_enqValid( T798 ),
       .io_deqValid( CU_24_io_deqValid ),
       .io_enqRdyOut( CU_24_io_enqRdyOut )
  );
  Switch_0 Switch(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       .io_inPort_4( CU_io_out ),
       .io_inPort_3( io_inData_0 ),
       //.io_inPort_2(  )
       .io_inPort_1( Switch_1_io_outPort_3 ),
       .io_inPort_0( Switch_6_io_outPort_2 ),
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       .io_outPort_4( Switch_io_outPort_4 ),
       .io_outPort_3( Switch_io_outPort_3 ),
       //.io_outPort_2(  )
       .io_outPort_1( Switch_io_outPort_1 ),
       .io_outPort_0( Switch_io_outPort_0 ),
       .io_deqValid( Switch_io_deqValid ),
       .io_enqRdy( Switch_io_enqRdy ),
       .io_deqRdy( T791 ),
       .io_enqValid( T784 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_io_outCUConfig ),
       .io_deqOR( Switch_1_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T783 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch.io_inPort_7 = {2{$random}};
    assign Switch.io_inPort_6 = {2{$random}};
    assign Switch.io_inPort_5 = {2{$random}};
    assign Switch.io_inPort_2 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_1(.clk(clk), .reset(reset),
       .io_inPort_7( CU_io_out ),
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       .io_inPort_4( CU_1_io_out ),
       .io_inPort_3( Switch_io_outPort_1 ),
       .io_inPort_2( io_inData_19 ),
       .io_inPort_1( Switch_2_io_outPort_3 ),
       .io_inPort_0( Switch_7_io_outPort_2 ),
       .io_outPort_7( Switch_1_io_outPort_7 ),
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       .io_outPort_4( Switch_1_io_outPort_4 ),
       .io_outPort_3( Switch_1_io_outPort_3 ),
       .io_outPort_2( Switch_1_io_outPort_2 ),
       .io_outPort_1( Switch_1_io_outPort_1 ),
       .io_outPort_0( Switch_1_io_outPort_0 ),
       .io_deqValid( Switch_1_io_deqValid ),
       .io_enqRdy( Switch_1_io_enqRdy ),
       .io_deqRdy( T774 ),
       .io_enqValid( T765 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_1_io_outCUConfig ),
       .io_deqOR( Switch_2_io_enqOR ),
       .io_enqOR( Switch_1_io_enqOR ),
       .io_deqRdyOut( T763 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_1.io_inPort_6 = {2{$random}};
    assign Switch_1.io_inPort_5 = {2{$random}};
// synthesis translate_on
`endif
  Switch_2 Switch_2(.clk(clk), .reset(reset),
       .io_inPort_7( CU_1_io_out ),
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       .io_inPort_4( CU_2_io_out ),
       .io_inPort_3( Switch_1_io_outPort_1 ),
       .io_inPort_2( io_inData_18 ),
       .io_inPort_1( Switch_3_io_outPort_3 ),
       .io_inPort_0( Switch_8_io_outPort_2 ),
       .io_outPort_7( Switch_2_io_outPort_7 ),
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       .io_outPort_4( Switch_2_io_outPort_4 ),
       .io_outPort_3( Switch_2_io_outPort_3 ),
       .io_outPort_2( Switch_2_io_outPort_2 ),
       .io_outPort_1( Switch_2_io_outPort_1 ),
       .io_outPort_0( Switch_2_io_outPort_0 ),
       .io_deqValid( Switch_2_io_deqValid ),
       .io_enqRdy( Switch_2_io_enqRdy ),
       .io_deqRdy( T754 ),
       .io_enqValid( T745 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_2_io_outCUConfig ),
       .io_deqOR( Switch_3_io_enqOR ),
       .io_enqOR( Switch_2_io_enqOR ),
       .io_deqRdyOut( T743 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_2.io_inPort_6 = {2{$random}};
    assign Switch_2.io_inPort_5 = {2{$random}};
// synthesis translate_on
`endif
  Switch_3 Switch_3(.clk(clk), .reset(reset),
       .io_inPort_7( CU_2_io_out ),
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       .io_inPort_4( CU_3_io_out ),
       .io_inPort_3( Switch_2_io_outPort_1 ),
       .io_inPort_2( io_inData_17 ),
       .io_inPort_1( Switch_4_io_outPort_3 ),
       .io_inPort_0( Switch_9_io_outPort_2 ),
       .io_outPort_7( Switch_3_io_outPort_7 ),
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       .io_outPort_4( Switch_3_io_outPort_4 ),
       .io_outPort_3( Switch_3_io_outPort_3 ),
       .io_outPort_2( Switch_3_io_outPort_2 ),
       .io_outPort_1( Switch_3_io_outPort_1 ),
       .io_outPort_0( Switch_3_io_outPort_0 ),
       .io_deqValid( Switch_3_io_deqValid ),
       .io_enqRdy( Switch_3_io_enqRdy ),
       .io_deqRdy( T734 ),
       .io_enqValid( T725 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_3_io_outCUConfig ),
       .io_deqOR( Switch_4_io_enqOR ),
       .io_enqOR( Switch_3_io_enqOR ),
       .io_deqRdyOut( T723 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_3.io_inPort_6 = {2{$random}};
    assign Switch_3.io_inPort_5 = {2{$random}};
// synthesis translate_on
`endif
  Switch_4 Switch_4(.clk(clk), .reset(reset),
       .io_inPort_7( CU_3_io_out ),
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       .io_inPort_4( CU_4_io_out ),
       .io_inPort_3( Switch_3_io_outPort_1 ),
       .io_inPort_2( io_inData_16 ),
       .io_inPort_1( Switch_5_io_outPort_3 ),
       .io_inPort_0( Switch_10_io_outPort_2 ),
       .io_outPort_7( Switch_4_io_outPort_7 ),
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       .io_outPort_4( Switch_4_io_outPort_4 ),
       .io_outPort_3( Switch_4_io_outPort_3 ),
       .io_outPort_2( Switch_4_io_outPort_2 ),
       .io_outPort_1( Switch_4_io_outPort_1 ),
       .io_outPort_0( Switch_4_io_outPort_0 ),
       .io_deqValid( Switch_4_io_deqValid ),
       .io_enqRdy( Switch_4_io_enqRdy ),
       .io_deqRdy( T714 ),
       .io_enqValid( T705 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_4_io_outCUConfig ),
       .io_deqOR( Switch_5_io_enqOR ),
       .io_enqOR( Switch_4_io_enqOR ),
       .io_deqRdyOut( T703 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_4.io_inPort_6 = {2{$random}};
    assign Switch_4.io_inPort_5 = {2{$random}};
// synthesis translate_on
`endif
  Switch_5 Switch_5(.clk(clk), .reset(reset),
       .io_inPort_7( CU_4_io_out ),
       //.io_inPort_6(  )
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_4_io_outPort_1 ),
       //.io_inPort_2(  )
       .io_inPort_1( io_inData_15 ),
       .io_inPort_0( Switch_11_io_outPort_2 ),
       .io_outPort_7( Switch_5_io_outPort_7 ),
       //.io_outPort_6(  )
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_5_io_outPort_3 ),
       //.io_outPort_2(  )
       .io_outPort_1( Switch_5_io_outPort_1 ),
       .io_outPort_0( Switch_5_io_outPort_0 ),
       .io_deqValid( Switch_5_io_deqValid ),
       .io_enqRdy( Switch_5_io_enqRdy ),
       .io_deqRdy( T696 ),
       .io_enqValid( T689 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_5_io_enqOR ),
       .io_deqRdyOut( T688 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_5.io_inPort_6 = {2{$random}};
    assign Switch_5.io_inPort_5 = {2{$random}};
    assign Switch_5.io_inPort_4 = {2{$random}};
    assign Switch_5.io_inPort_2 = {2{$random}};
// synthesis translate_on
`endif
  Switch_0 Switch_6(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       .io_inPort_5( CU_io_out ),
       .io_inPort_4( CU_5_io_out ),
       .io_inPort_3( io_inData_1 ),
       .io_inPort_2( Switch_io_outPort_0 ),
       .io_inPort_1( Switch_7_io_outPort_3 ),
       .io_inPort_0( Switch_12_io_outPort_2 ),
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       .io_outPort_5( Switch_6_io_outPort_5 ),
       .io_outPort_4( Switch_6_io_outPort_4 ),
       .io_outPort_3( Switch_6_io_outPort_3 ),
       .io_outPort_2( Switch_6_io_outPort_2 ),
       .io_outPort_1( Switch_6_io_outPort_1 ),
       .io_outPort_0( Switch_6_io_outPort_0 ),
       .io_deqValid( Switch_6_io_deqValid ),
       .io_enqRdy( Switch_6_io_enqRdy ),
       .io_deqRdy( T679 ),
       .io_enqValid( T670 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_6_io_outCUConfig ),
       .io_deqOR( Switch_7_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T668 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_6.io_inPort_7 = {2{$random}};
    assign Switch_6.io_inPort_6 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_7(.clk(clk), .reset(reset),
       .io_inPort_7( CU_5_io_out ),
       .io_inPort_6( CU_io_out ),
       .io_inPort_5( CU_1_io_out ),
       .io_inPort_4( CU_6_io_out ),
       .io_inPort_3( Switch_6_io_outPort_1 ),
       .io_inPort_2( Switch_1_io_outPort_0 ),
       .io_inPort_1( Switch_8_io_outPort_3 ),
       .io_inPort_0( Switch_13_io_outPort_2 ),
       .io_outPort_7( Switch_7_io_outPort_7 ),
       .io_outPort_6( Switch_7_io_outPort_6 ),
       .io_outPort_5( Switch_7_io_outPort_5 ),
       .io_outPort_4( Switch_7_io_outPort_4 ),
       .io_outPort_3( Switch_7_io_outPort_3 ),
       .io_outPort_2( Switch_7_io_outPort_2 ),
       .io_outPort_1( Switch_7_io_outPort_1 ),
       .io_outPort_0( Switch_7_io_outPort_0 ),
       .io_deqValid( Switch_7_io_deqValid ),
       .io_enqRdy( Switch_7_io_enqRdy ),
       .io_deqRdy( T657 ),
       .io_enqValid( T646 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_7_io_outCUConfig ),
       .io_deqOR( Switch_8_io_enqOR ),
       .io_enqOR( Switch_7_io_enqOR ),
       .io_deqRdyOut( T643 )
  );
  Switch_2 Switch_8(.clk(clk), .reset(reset),
       .io_inPort_7( CU_6_io_out ),
       .io_inPort_6( CU_1_io_out ),
       .io_inPort_5( CU_2_io_out ),
       .io_inPort_4( CU_7_io_out ),
       .io_inPort_3( Switch_7_io_outPort_1 ),
       .io_inPort_2( Switch_2_io_outPort_0 ),
       .io_inPort_1( Switch_9_io_outPort_3 ),
       .io_inPort_0( Switch_14_io_outPort_2 ),
       .io_outPort_7( Switch_8_io_outPort_7 ),
       .io_outPort_6( Switch_8_io_outPort_6 ),
       .io_outPort_5( Switch_8_io_outPort_5 ),
       .io_outPort_4( Switch_8_io_outPort_4 ),
       .io_outPort_3( Switch_8_io_outPort_3 ),
       .io_outPort_2( Switch_8_io_outPort_2 ),
       .io_outPort_1( Switch_8_io_outPort_1 ),
       .io_outPort_0( Switch_8_io_outPort_0 ),
       .io_deqValid( Switch_8_io_deqValid ),
       .io_enqRdy( Switch_8_io_enqRdy ),
       .io_deqRdy( T632 ),
       .io_enqValid( T621 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_8_io_outCUConfig ),
       .io_deqOR( Switch_9_io_enqOR ),
       .io_enqOR( Switch_8_io_enqOR ),
       .io_deqRdyOut( T618 )
  );
  Switch_3 Switch_9(.clk(clk), .reset(reset),
       .io_inPort_7( CU_7_io_out ),
       .io_inPort_6( CU_2_io_out ),
       .io_inPort_5( CU_3_io_out ),
       .io_inPort_4( CU_8_io_out ),
       .io_inPort_3( Switch_8_io_outPort_1 ),
       .io_inPort_2( Switch_3_io_outPort_0 ),
       .io_inPort_1( Switch_10_io_outPort_3 ),
       .io_inPort_0( Switch_15_io_outPort_2 ),
       .io_outPort_7( Switch_9_io_outPort_7 ),
       .io_outPort_6( Switch_9_io_outPort_6 ),
       .io_outPort_5( Switch_9_io_outPort_5 ),
       .io_outPort_4( Switch_9_io_outPort_4 ),
       .io_outPort_3( Switch_9_io_outPort_3 ),
       .io_outPort_2( Switch_9_io_outPort_2 ),
       .io_outPort_1( Switch_9_io_outPort_1 ),
       .io_outPort_0( Switch_9_io_outPort_0 ),
       .io_deqValid( Switch_9_io_deqValid ),
       .io_enqRdy( Switch_9_io_enqRdy ),
       .io_deqRdy( T607 ),
       .io_enqValid( T596 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_9_io_outCUConfig ),
       .io_deqOR( Switch_10_io_enqOR ),
       .io_enqOR( Switch_9_io_enqOR ),
       .io_deqRdyOut( T593 )
  );
  Switch_4 Switch_10(.clk(clk), .reset(reset),
       .io_inPort_7( CU_8_io_out ),
       .io_inPort_6( CU_3_io_out ),
       .io_inPort_5( CU_4_io_out ),
       .io_inPort_4( CU_9_io_out ),
       .io_inPort_3( Switch_9_io_outPort_1 ),
       .io_inPort_2( Switch_4_io_outPort_0 ),
       .io_inPort_1( Switch_11_io_outPort_3 ),
       .io_inPort_0( Switch_16_io_outPort_2 ),
       .io_outPort_7( Switch_10_io_outPort_7 ),
       .io_outPort_6( Switch_10_io_outPort_6 ),
       .io_outPort_5( Switch_10_io_outPort_5 ),
       .io_outPort_4( Switch_10_io_outPort_4 ),
       .io_outPort_3( Switch_10_io_outPort_3 ),
       .io_outPort_2( Switch_10_io_outPort_2 ),
       .io_outPort_1( Switch_10_io_outPort_1 ),
       .io_outPort_0( Switch_10_io_outPort_0 ),
       .io_deqValid( Switch_10_io_deqValid ),
       .io_enqRdy( Switch_10_io_enqRdy ),
       .io_deqRdy( T582 ),
       .io_enqValid( T571 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_10_io_outCUConfig ),
       .io_deqOR( Switch_11_io_enqOR ),
       .io_enqOR( Switch_10_io_enqOR ),
       .io_deqRdyOut( T568 )
  );
  Switch_5 Switch_11(.clk(clk), .reset(reset),
       .io_inPort_7( CU_9_io_out ),
       .io_inPort_6( CU_4_io_out ),
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_10_io_outPort_1 ),
       .io_inPort_2( Switch_5_io_outPort_0 ),
       .io_inPort_1( io_inData_14 ),
       .io_inPort_0( Switch_17_io_outPort_2 ),
       .io_outPort_7( Switch_11_io_outPort_7 ),
       .io_outPort_6( Switch_11_io_outPort_6 ),
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_11_io_outPort_3 ),
       .io_outPort_2( Switch_11_io_outPort_2 ),
       .io_outPort_1( Switch_11_io_outPort_1 ),
       .io_outPort_0( Switch_11_io_outPort_0 ),
       .io_deqValid( Switch_11_io_deqValid ),
       .io_enqRdy( Switch_11_io_enqRdy ),
       .io_deqRdy( T559 ),
       .io_enqValid( T550 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_11_io_enqOR ),
       .io_deqRdyOut( T548 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_11.io_inPort_5 = {2{$random}};
    assign Switch_11.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_0 Switch_12(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       .io_inPort_5( CU_5_io_out ),
       .io_inPort_4( CU_10_io_out ),
       .io_inPort_3( io_inData_2 ),
       .io_inPort_2( Switch_6_io_outPort_0 ),
       .io_inPort_1( Switch_13_io_outPort_3 ),
       .io_inPort_0( Switch_18_io_outPort_2 ),
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       .io_outPort_5( Switch_12_io_outPort_5 ),
       .io_outPort_4( Switch_12_io_outPort_4 ),
       .io_outPort_3( Switch_12_io_outPort_3 ),
       .io_outPort_2( Switch_12_io_outPort_2 ),
       .io_outPort_1( Switch_12_io_outPort_1 ),
       .io_outPort_0( Switch_12_io_outPort_0 ),
       .io_deqValid( Switch_12_io_deqValid ),
       .io_enqRdy( Switch_12_io_enqRdy ),
       .io_deqRdy( T539 ),
       .io_enqValid( T530 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_12_io_outCUConfig ),
       .io_deqOR( Switch_13_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T528 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_12.io_inPort_7 = {2{$random}};
    assign Switch_12.io_inPort_6 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_13(.clk(clk), .reset(reset),
       .io_inPort_7( CU_10_io_out ),
       .io_inPort_6( CU_5_io_out ),
       .io_inPort_5( CU_6_io_out ),
       .io_inPort_4( CU_11_io_out ),
       .io_inPort_3( Switch_12_io_outPort_1 ),
       .io_inPort_2( Switch_7_io_outPort_0 ),
       .io_inPort_1( Switch_14_io_outPort_3 ),
       .io_inPort_0( Switch_19_io_outPort_2 ),
       .io_outPort_7( Switch_13_io_outPort_7 ),
       .io_outPort_6( Switch_13_io_outPort_6 ),
       .io_outPort_5( Switch_13_io_outPort_5 ),
       .io_outPort_4( Switch_13_io_outPort_4 ),
       .io_outPort_3( Switch_13_io_outPort_3 ),
       .io_outPort_2( Switch_13_io_outPort_2 ),
       .io_outPort_1( Switch_13_io_outPort_1 ),
       .io_outPort_0( Switch_13_io_outPort_0 ),
       .io_deqValid( Switch_13_io_deqValid ),
       .io_enqRdy( Switch_13_io_enqRdy ),
       .io_deqRdy( T517 ),
       .io_enqValid( T506 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_13_io_outCUConfig ),
       .io_deqOR( Switch_14_io_enqOR ),
       .io_enqOR( Switch_13_io_enqOR ),
       .io_deqRdyOut( T503 )
  );
  Switch_2 Switch_14(.clk(clk), .reset(reset),
       .io_inPort_7( CU_11_io_out ),
       .io_inPort_6( CU_6_io_out ),
       .io_inPort_5( CU_7_io_out ),
       .io_inPort_4( CU_12_io_out ),
       .io_inPort_3( Switch_13_io_outPort_1 ),
       .io_inPort_2( Switch_8_io_outPort_0 ),
       .io_inPort_1( Switch_15_io_outPort_3 ),
       .io_inPort_0( Switch_20_io_outPort_2 ),
       .io_outPort_7( Switch_14_io_outPort_7 ),
       .io_outPort_6( Switch_14_io_outPort_6 ),
       .io_outPort_5( Switch_14_io_outPort_5 ),
       .io_outPort_4( Switch_14_io_outPort_4 ),
       .io_outPort_3( Switch_14_io_outPort_3 ),
       .io_outPort_2( Switch_14_io_outPort_2 ),
       .io_outPort_1( Switch_14_io_outPort_1 ),
       .io_outPort_0( Switch_14_io_outPort_0 ),
       .io_deqValid( Switch_14_io_deqValid ),
       .io_enqRdy( Switch_14_io_enqRdy ),
       .io_deqRdy( T492 ),
       .io_enqValid( T481 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_14_io_outCUConfig ),
       .io_deqOR( Switch_15_io_enqOR ),
       .io_enqOR( Switch_14_io_enqOR ),
       .io_deqRdyOut( T478 )
  );
  Switch_3 Switch_15(.clk(clk), .reset(reset),
       .io_inPort_7( CU_12_io_out ),
       .io_inPort_6( CU_7_io_out ),
       .io_inPort_5( CU_8_io_out ),
       .io_inPort_4( CU_13_io_out ),
       .io_inPort_3( Switch_14_io_outPort_1 ),
       .io_inPort_2( Switch_9_io_outPort_0 ),
       .io_inPort_1( Switch_16_io_outPort_3 ),
       .io_inPort_0( Switch_21_io_outPort_2 ),
       .io_outPort_7( Switch_15_io_outPort_7 ),
       .io_outPort_6( Switch_15_io_outPort_6 ),
       .io_outPort_5( Switch_15_io_outPort_5 ),
       .io_outPort_4( Switch_15_io_outPort_4 ),
       .io_outPort_3( Switch_15_io_outPort_3 ),
       .io_outPort_2( Switch_15_io_outPort_2 ),
       .io_outPort_1( Switch_15_io_outPort_1 ),
       .io_outPort_0( Switch_15_io_outPort_0 ),
       .io_deqValid( Switch_15_io_deqValid ),
       .io_enqRdy( Switch_15_io_enqRdy ),
       .io_deqRdy( T467 ),
       .io_enqValid( T456 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_15_io_outCUConfig ),
       .io_deqOR( Switch_16_io_enqOR ),
       .io_enqOR( Switch_15_io_enqOR ),
       .io_deqRdyOut( T453 )
  );
  Switch_4 Switch_16(.clk(clk), .reset(reset),
       .io_inPort_7( CU_13_io_out ),
       .io_inPort_6( CU_8_io_out ),
       .io_inPort_5( CU_9_io_out ),
       .io_inPort_4( CU_14_io_out ),
       .io_inPort_3( Switch_15_io_outPort_1 ),
       .io_inPort_2( Switch_10_io_outPort_0 ),
       .io_inPort_1( Switch_17_io_outPort_3 ),
       .io_inPort_0( Switch_22_io_outPort_2 ),
       .io_outPort_7( Switch_16_io_outPort_7 ),
       .io_outPort_6( Switch_16_io_outPort_6 ),
       .io_outPort_5( Switch_16_io_outPort_5 ),
       .io_outPort_4( Switch_16_io_outPort_4 ),
       .io_outPort_3( Switch_16_io_outPort_3 ),
       .io_outPort_2( Switch_16_io_outPort_2 ),
       .io_outPort_1( Switch_16_io_outPort_1 ),
       .io_outPort_0( Switch_16_io_outPort_0 ),
       .io_deqValid( Switch_16_io_deqValid ),
       .io_enqRdy( Switch_16_io_enqRdy ),
       .io_deqRdy( T442 ),
       .io_enqValid( T431 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_16_io_outCUConfig ),
       .io_deqOR( Switch_17_io_enqOR ),
       .io_enqOR( Switch_16_io_enqOR ),
       .io_deqRdyOut( T428 )
  );
  Switch_5 Switch_17(.clk(clk), .reset(reset),
       .io_inPort_7( CU_14_io_out ),
       .io_inPort_6( CU_9_io_out ),
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_16_io_outPort_1 ),
       .io_inPort_2( Switch_11_io_outPort_0 ),
       .io_inPort_1( io_inData_13 ),
       .io_inPort_0( Switch_23_io_outPort_2 ),
       .io_outPort_7( Switch_17_io_outPort_7 ),
       .io_outPort_6( Switch_17_io_outPort_6 ),
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_17_io_outPort_3 ),
       .io_outPort_2( Switch_17_io_outPort_2 ),
       .io_outPort_1( Switch_17_io_outPort_1 ),
       .io_outPort_0( Switch_17_io_outPort_0 ),
       .io_deqValid( Switch_17_io_deqValid ),
       .io_enqRdy( Switch_17_io_enqRdy ),
       .io_deqRdy( T419 ),
       .io_enqValid( T410 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_17_io_enqOR ),
       .io_deqRdyOut( T408 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_17.io_inPort_5 = {2{$random}};
    assign Switch_17.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_0 Switch_18(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       .io_inPort_5( CU_10_io_out ),
       .io_inPort_4( CU_15_io_out ),
       .io_inPort_3( io_inData_3 ),
       .io_inPort_2( Switch_12_io_outPort_0 ),
       .io_inPort_1( Switch_19_io_outPort_3 ),
       .io_inPort_0( Switch_24_io_outPort_2 ),
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       .io_outPort_5( Switch_18_io_outPort_5 ),
       .io_outPort_4( Switch_18_io_outPort_4 ),
       .io_outPort_3( Switch_18_io_outPort_3 ),
       .io_outPort_2( Switch_18_io_outPort_2 ),
       .io_outPort_1( Switch_18_io_outPort_1 ),
       .io_outPort_0( Switch_18_io_outPort_0 ),
       .io_deqValid( Switch_18_io_deqValid ),
       .io_enqRdy( Switch_18_io_enqRdy ),
       .io_deqRdy( T399 ),
       .io_enqValid( T390 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_18_io_outCUConfig ),
       .io_deqOR( Switch_19_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T388 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_18.io_inPort_7 = {2{$random}};
    assign Switch_18.io_inPort_6 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_19(.clk(clk), .reset(reset),
       .io_inPort_7( CU_15_io_out ),
       .io_inPort_6( CU_10_io_out ),
       .io_inPort_5( CU_11_io_out ),
       .io_inPort_4( CU_16_io_out ),
       .io_inPort_3( Switch_18_io_outPort_1 ),
       .io_inPort_2( Switch_13_io_outPort_0 ),
       .io_inPort_1( Switch_20_io_outPort_3 ),
       .io_inPort_0( Switch_25_io_outPort_2 ),
       .io_outPort_7( Switch_19_io_outPort_7 ),
       .io_outPort_6( Switch_19_io_outPort_6 ),
       .io_outPort_5( Switch_19_io_outPort_5 ),
       .io_outPort_4( Switch_19_io_outPort_4 ),
       .io_outPort_3( Switch_19_io_outPort_3 ),
       .io_outPort_2( Switch_19_io_outPort_2 ),
       .io_outPort_1( Switch_19_io_outPort_1 ),
       .io_outPort_0( Switch_19_io_outPort_0 ),
       .io_deqValid( Switch_19_io_deqValid ),
       .io_enqRdy( Switch_19_io_enqRdy ),
       .io_deqRdy( T377 ),
       .io_enqValid( T366 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_19_io_outCUConfig ),
       .io_deqOR( Switch_20_io_enqOR ),
       .io_enqOR( Switch_19_io_enqOR ),
       .io_deqRdyOut( T363 )
  );
  Switch_2 Switch_20(.clk(clk), .reset(reset),
       .io_inPort_7( CU_16_io_out ),
       .io_inPort_6( CU_11_io_out ),
       .io_inPort_5( CU_12_io_out ),
       .io_inPort_4( CU_17_io_out ),
       .io_inPort_3( Switch_19_io_outPort_1 ),
       .io_inPort_2( Switch_14_io_outPort_0 ),
       .io_inPort_1( Switch_21_io_outPort_3 ),
       .io_inPort_0( Switch_26_io_outPort_2 ),
       .io_outPort_7( Switch_20_io_outPort_7 ),
       .io_outPort_6( Switch_20_io_outPort_6 ),
       .io_outPort_5( Switch_20_io_outPort_5 ),
       .io_outPort_4( Switch_20_io_outPort_4 ),
       .io_outPort_3( Switch_20_io_outPort_3 ),
       .io_outPort_2( Switch_20_io_outPort_2 ),
       .io_outPort_1( Switch_20_io_outPort_1 ),
       .io_outPort_0( Switch_20_io_outPort_0 ),
       .io_deqValid( Switch_20_io_deqValid ),
       .io_enqRdy( Switch_20_io_enqRdy ),
       .io_deqRdy( T352 ),
       .io_enqValid( T341 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_20_io_outCUConfig ),
       .io_deqOR( Switch_21_io_enqOR ),
       .io_enqOR( Switch_20_io_enqOR ),
       .io_deqRdyOut( T338 )
  );
  Switch_3 Switch_21(.clk(clk), .reset(reset),
       .io_inPort_7( CU_17_io_out ),
       .io_inPort_6( CU_12_io_out ),
       .io_inPort_5( CU_13_io_out ),
       .io_inPort_4( CU_18_io_out ),
       .io_inPort_3( Switch_20_io_outPort_1 ),
       .io_inPort_2( Switch_15_io_outPort_0 ),
       .io_inPort_1( Switch_22_io_outPort_3 ),
       .io_inPort_0( Switch_27_io_outPort_2 ),
       .io_outPort_7( Switch_21_io_outPort_7 ),
       .io_outPort_6( Switch_21_io_outPort_6 ),
       .io_outPort_5( Switch_21_io_outPort_5 ),
       .io_outPort_4( Switch_21_io_outPort_4 ),
       .io_outPort_3( Switch_21_io_outPort_3 ),
       .io_outPort_2( Switch_21_io_outPort_2 ),
       .io_outPort_1( Switch_21_io_outPort_1 ),
       .io_outPort_0( Switch_21_io_outPort_0 ),
       .io_deqValid( Switch_21_io_deqValid ),
       .io_enqRdy( Switch_21_io_enqRdy ),
       .io_deqRdy( T327 ),
       .io_enqValid( T316 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_21_io_outCUConfig ),
       .io_deqOR( Switch_22_io_enqOR ),
       .io_enqOR( Switch_21_io_enqOR ),
       .io_deqRdyOut( T313 )
  );
  Switch_4 Switch_22(.clk(clk), .reset(reset),
       .io_inPort_7( CU_18_io_out ),
       .io_inPort_6( CU_13_io_out ),
       .io_inPort_5( CU_14_io_out ),
       .io_inPort_4( CU_19_io_out ),
       .io_inPort_3( Switch_21_io_outPort_1 ),
       .io_inPort_2( Switch_16_io_outPort_0 ),
       .io_inPort_1( Switch_23_io_outPort_3 ),
       .io_inPort_0( Switch_28_io_outPort_2 ),
       .io_outPort_7( Switch_22_io_outPort_7 ),
       .io_outPort_6( Switch_22_io_outPort_6 ),
       .io_outPort_5( Switch_22_io_outPort_5 ),
       .io_outPort_4( Switch_22_io_outPort_4 ),
       .io_outPort_3( Switch_22_io_outPort_3 ),
       .io_outPort_2( Switch_22_io_outPort_2 ),
       .io_outPort_1( Switch_22_io_outPort_1 ),
       .io_outPort_0( Switch_22_io_outPort_0 ),
       .io_deqValid( Switch_22_io_deqValid ),
       .io_enqRdy( Switch_22_io_enqRdy ),
       .io_deqRdy( T302 ),
       .io_enqValid( T291 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_22_io_outCUConfig ),
       .io_deqOR( Switch_23_io_enqOR ),
       .io_enqOR( Switch_22_io_enqOR ),
       .io_deqRdyOut( T288 )
  );
  Switch_5 Switch_23(.clk(clk), .reset(reset),
       .io_inPort_7( CU_19_io_out ),
       .io_inPort_6( CU_14_io_out ),
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_22_io_outPort_1 ),
       .io_inPort_2( Switch_17_io_outPort_0 ),
       .io_inPort_1( io_inData_12 ),
       .io_inPort_0( Switch_29_io_outPort_2 ),
       .io_outPort_7( Switch_23_io_outPort_7 ),
       .io_outPort_6( Switch_23_io_outPort_6 ),
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_23_io_outPort_3 ),
       .io_outPort_2( Switch_23_io_outPort_2 ),
       .io_outPort_1( Switch_23_io_outPort_1 ),
       .io_outPort_0( Switch_23_io_outPort_0 ),
       .io_deqValid( Switch_23_io_deqValid ),
       .io_enqRdy( Switch_23_io_enqRdy ),
       .io_deqRdy( T279 ),
       .io_enqValid( T270 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_23_io_enqOR ),
       .io_deqRdyOut( T268 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_23.io_inPort_5 = {2{$random}};
    assign Switch_23.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_0 Switch_24(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       .io_inPort_5( CU_15_io_out ),
       .io_inPort_4( CU_20_io_out ),
       .io_inPort_3( io_inData_4 ),
       .io_inPort_2( Switch_18_io_outPort_0 ),
       .io_inPort_1( Switch_25_io_outPort_3 ),
       .io_inPort_0( Switch_30_io_outPort_2 ),
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       .io_outPort_5( Switch_24_io_outPort_5 ),
       .io_outPort_4( Switch_24_io_outPort_4 ),
       .io_outPort_3( Switch_24_io_outPort_3 ),
       .io_outPort_2( Switch_24_io_outPort_2 ),
       .io_outPort_1( Switch_24_io_outPort_1 ),
       .io_outPort_0( Switch_24_io_outPort_0 ),
       .io_deqValid( Switch_24_io_deqValid ),
       .io_enqRdy( Switch_24_io_enqRdy ),
       .io_deqRdy( T259 ),
       .io_enqValid( T250 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_24_io_outCUConfig ),
       .io_deqOR( Switch_25_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T248 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_24.io_inPort_7 = {2{$random}};
    assign Switch_24.io_inPort_6 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_25(.clk(clk), .reset(reset),
       .io_inPort_7( CU_20_io_out ),
       .io_inPort_6( CU_15_io_out ),
       .io_inPort_5( CU_16_io_out ),
       .io_inPort_4( CU_21_io_out ),
       .io_inPort_3( Switch_24_io_outPort_1 ),
       .io_inPort_2( Switch_19_io_outPort_0 ),
       .io_inPort_1( Switch_26_io_outPort_3 ),
       .io_inPort_0( Switch_31_io_outPort_2 ),
       .io_outPort_7( Switch_25_io_outPort_7 ),
       .io_outPort_6( Switch_25_io_outPort_6 ),
       .io_outPort_5( Switch_25_io_outPort_5 ),
       .io_outPort_4( Switch_25_io_outPort_4 ),
       .io_outPort_3( Switch_25_io_outPort_3 ),
       .io_outPort_2( Switch_25_io_outPort_2 ),
       .io_outPort_1( Switch_25_io_outPort_1 ),
       .io_outPort_0( Switch_25_io_outPort_0 ),
       .io_deqValid( Switch_25_io_deqValid ),
       .io_enqRdy( Switch_25_io_enqRdy ),
       .io_deqRdy( T237 ),
       .io_enqValid( T226 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_25_io_outCUConfig ),
       .io_deqOR( Switch_26_io_enqOR ),
       .io_enqOR( Switch_25_io_enqOR ),
       .io_deqRdyOut( T223 )
  );
  Switch_2 Switch_26(.clk(clk), .reset(reset),
       .io_inPort_7( CU_21_io_out ),
       .io_inPort_6( CU_16_io_out ),
       .io_inPort_5( CU_17_io_out ),
       .io_inPort_4( CU_22_io_out ),
       .io_inPort_3( Switch_25_io_outPort_1 ),
       .io_inPort_2( Switch_20_io_outPort_0 ),
       .io_inPort_1( Switch_27_io_outPort_3 ),
       .io_inPort_0( Switch_32_io_outPort_2 ),
       .io_outPort_7( Switch_26_io_outPort_7 ),
       .io_outPort_6( Switch_26_io_outPort_6 ),
       .io_outPort_5( Switch_26_io_outPort_5 ),
       .io_outPort_4( Switch_26_io_outPort_4 ),
       .io_outPort_3( Switch_26_io_outPort_3 ),
       .io_outPort_2( Switch_26_io_outPort_2 ),
       .io_outPort_1( Switch_26_io_outPort_1 ),
       .io_outPort_0( Switch_26_io_outPort_0 ),
       .io_deqValid( Switch_26_io_deqValid ),
       .io_enqRdy( Switch_26_io_enqRdy ),
       .io_deqRdy( T212 ),
       .io_enqValid( T201 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_26_io_outCUConfig ),
       .io_deqOR( Switch_27_io_enqOR ),
       .io_enqOR( Switch_26_io_enqOR ),
       .io_deqRdyOut( T198 )
  );
  Switch_3 Switch_27(.clk(clk), .reset(reset),
       .io_inPort_7( CU_22_io_out ),
       .io_inPort_6( CU_17_io_out ),
       .io_inPort_5( CU_18_io_out ),
       .io_inPort_4( CU_23_io_out ),
       .io_inPort_3( Switch_26_io_outPort_1 ),
       .io_inPort_2( Switch_21_io_outPort_0 ),
       .io_inPort_1( Switch_28_io_outPort_3 ),
       .io_inPort_0( Switch_33_io_outPort_2 ),
       .io_outPort_7( Switch_27_io_outPort_7 ),
       .io_outPort_6( Switch_27_io_outPort_6 ),
       .io_outPort_5( Switch_27_io_outPort_5 ),
       .io_outPort_4( Switch_27_io_outPort_4 ),
       .io_outPort_3( Switch_27_io_outPort_3 ),
       .io_outPort_2( Switch_27_io_outPort_2 ),
       .io_outPort_1( Switch_27_io_outPort_1 ),
       .io_outPort_0( Switch_27_io_outPort_0 ),
       .io_deqValid( Switch_27_io_deqValid ),
       .io_enqRdy( Switch_27_io_enqRdy ),
       .io_deqRdy( T187 ),
       .io_enqValid( T176 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_27_io_outCUConfig ),
       .io_deqOR( Switch_28_io_enqOR ),
       .io_enqOR( Switch_27_io_enqOR ),
       .io_deqRdyOut( T173 )
  );
  Switch_4 Switch_28(.clk(clk), .reset(reset),
       .io_inPort_7( CU_23_io_out ),
       .io_inPort_6( CU_18_io_out ),
       .io_inPort_5( CU_19_io_out ),
       .io_inPort_4( CU_24_io_out ),
       .io_inPort_3( Switch_27_io_outPort_1 ),
       .io_inPort_2( Switch_22_io_outPort_0 ),
       .io_inPort_1( Switch_29_io_outPort_3 ),
       .io_inPort_0( Switch_34_io_outPort_2 ),
       .io_outPort_7( Switch_28_io_outPort_7 ),
       .io_outPort_6( Switch_28_io_outPort_6 ),
       .io_outPort_5( Switch_28_io_outPort_5 ),
       .io_outPort_4( Switch_28_io_outPort_4 ),
       .io_outPort_3( Switch_28_io_outPort_3 ),
       .io_outPort_2( Switch_28_io_outPort_2 ),
       .io_outPort_1( Switch_28_io_outPort_1 ),
       .io_outPort_0( Switch_28_io_outPort_0 ),
       .io_deqValid( Switch_28_io_deqValid ),
       .io_enqRdy( Switch_28_io_enqRdy ),
       .io_deqRdy( T162 ),
       .io_enqValid( T151 ),
       //.io_outConfigData(  )
       .io_outCUConfig( Switch_28_io_outCUConfig ),
       .io_deqOR( Switch_29_io_enqOR ),
       .io_enqOR( Switch_28_io_enqOR ),
       .io_deqRdyOut( T148 )
  );
  Switch_5 Switch_29(.clk(clk), .reset(reset),
       .io_inPort_7( CU_24_io_out ),
       .io_inPort_6( CU_19_io_out ),
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_28_io_outPort_1 ),
       .io_inPort_2( Switch_23_io_outPort_0 ),
       .io_inPort_1( io_inData_11 ),
       .io_inPort_0( Switch_35_io_outPort_2 ),
       .io_outPort_7( Switch_29_io_outPort_7 ),
       .io_outPort_6( Switch_29_io_outPort_6 ),
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_29_io_outPort_3 ),
       .io_outPort_2( Switch_29_io_outPort_2 ),
       .io_outPort_1( Switch_29_io_outPort_1 ),
       .io_outPort_0( Switch_29_io_outPort_0 ),
       .io_deqValid( Switch_29_io_deqValid ),
       .io_enqRdy( Switch_29_io_enqRdy ),
       .io_deqRdy( T139 ),
       .io_enqValid( T130 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_29_io_enqOR ),
       .io_deqRdyOut( T128 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_29.io_inPort_5 = {2{$random}};
    assign Switch_29.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_0 Switch_30(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       //.io_inPort_6(  )
       .io_inPort_5( CU_20_io_out ),
       //.io_inPort_4(  )
       .io_inPort_3( io_inData_5 ),
       .io_inPort_2( Switch_24_io_outPort_0 ),
       .io_inPort_1( Switch_31_io_outPort_3 ),
       //.io_inPort_0(  )
       //.io_outPort_7(  )
       //.io_outPort_6(  )
       .io_outPort_5( Switch_30_io_outPort_5 ),
       //.io_outPort_4(  )
       .io_outPort_3( Switch_30_io_outPort_3 ),
       .io_outPort_2( Switch_30_io_outPort_2 ),
       .io_outPort_1( Switch_30_io_outPort_1 ),
       //.io_outPort_0(  )
       .io_deqValid( Switch_30_io_deqValid ),
       .io_enqRdy( Switch_30_io_enqRdy ),
       .io_deqRdy( T120 ),
       .io_enqValid( T112 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( Switch_31_io_enqOR ),
       //.io_enqOR(  )
       .io_deqRdyOut( T110 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_30.io_inPort_7 = {2{$random}};
    assign Switch_30.io_inPort_6 = {2{$random}};
    assign Switch_30.io_inPort_4 = {2{$random}};
    assign Switch_30.io_inPort_0 = {2{$random}};
// synthesis translate_on
`endif
  Switch_1 Switch_31(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       .io_inPort_6( CU_20_io_out ),
       .io_inPort_5( CU_21_io_out ),
       //.io_inPort_4(  )
       .io_inPort_3( Switch_30_io_outPort_1 ),
       .io_inPort_2( Switch_25_io_outPort_0 ),
       .io_inPort_1( Switch_32_io_outPort_3 ),
       .io_inPort_0( io_inData_6 ),
       //.io_outPort_7(  )
       .io_outPort_6( Switch_31_io_outPort_6 ),
       .io_outPort_5( Switch_31_io_outPort_5 ),
       //.io_outPort_4(  )
       .io_outPort_3( Switch_31_io_outPort_3 ),
       .io_outPort_2( Switch_31_io_outPort_2 ),
       .io_outPort_1( Switch_31_io_outPort_1 ),
       .io_outPort_0( Switch_31_io_outPort_0 ),
       .io_deqValid( Switch_31_io_deqValid ),
       .io_enqRdy( Switch_31_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( T90 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( Switch_32_io_enqOR ),
       .io_enqOR( Switch_31_io_enqOR ),
       .io_deqRdyOut( T87 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_31.io_inPort_7 = {2{$random}};
    assign Switch_31.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_2 Switch_32(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       .io_inPort_6( CU_21_io_out ),
       .io_inPort_5( CU_22_io_out ),
       //.io_inPort_4(  )
       .io_inPort_3( Switch_31_io_outPort_1 ),
       .io_inPort_2( Switch_26_io_outPort_0 ),
       .io_inPort_1( Switch_33_io_outPort_3 ),
       .io_inPort_0( io_inData_7 ),
       //.io_outPort_7(  )
       .io_outPort_6( Switch_32_io_outPort_6 ),
       .io_outPort_5( Switch_32_io_outPort_5 ),
       //.io_outPort_4(  )
       .io_outPort_3( Switch_32_io_outPort_3 ),
       .io_outPort_2( Switch_32_io_outPort_2 ),
       .io_outPort_1( Switch_32_io_outPort_1 ),
       .io_outPort_0( Switch_32_io_outPort_0 ),
       .io_deqValid( Switch_32_io_deqValid ),
       .io_enqRdy( Switch_32_io_enqRdy ),
       .io_deqRdy( T77 ),
       .io_enqValid( T67 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( Switch_33_io_enqOR ),
       .io_enqOR( Switch_32_io_enqOR ),
       .io_deqRdyOut( T64 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_32.io_inPort_7 = {2{$random}};
    assign Switch_32.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_3 Switch_33(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       .io_inPort_6( CU_22_io_out ),
       .io_inPort_5( CU_23_io_out ),
       //.io_inPort_4(  )
       .io_inPort_3( Switch_32_io_outPort_1 ),
       .io_inPort_2( Switch_27_io_outPort_0 ),
       .io_inPort_1( Switch_34_io_outPort_3 ),
       .io_inPort_0( io_inData_8 ),
       //.io_outPort_7(  )
       .io_outPort_6( Switch_33_io_outPort_6 ),
       .io_outPort_5( Switch_33_io_outPort_5 ),
       //.io_outPort_4(  )
       .io_outPort_3( Switch_33_io_outPort_3 ),
       .io_outPort_2( Switch_33_io_outPort_2 ),
       .io_outPort_1( Switch_33_io_outPort_1 ),
       .io_outPort_0( Switch_33_io_outPort_0 ),
       .io_deqValid( Switch_33_io_deqValid ),
       .io_enqRdy( Switch_33_io_enqRdy ),
       .io_deqRdy( T54 ),
       .io_enqValid( T44 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( Switch_34_io_enqOR ),
       .io_enqOR( Switch_33_io_enqOR ),
       .io_deqRdyOut( T41 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_33.io_inPort_7 = {2{$random}};
    assign Switch_33.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_4 Switch_34(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       .io_inPort_6( CU_23_io_out ),
       .io_inPort_5( CU_24_io_out ),
       //.io_inPort_4(  )
       .io_inPort_3( Switch_33_io_outPort_1 ),
       .io_inPort_2( Switch_28_io_outPort_0 ),
       .io_inPort_1( Switch_35_io_outPort_3 ),
       .io_inPort_0( io_inData_9 ),
       //.io_outPort_7(  )
       .io_outPort_6( Switch_34_io_outPort_6 ),
       .io_outPort_5( Switch_34_io_outPort_5 ),
       //.io_outPort_4(  )
       .io_outPort_3( Switch_34_io_outPort_3 ),
       .io_outPort_2( Switch_34_io_outPort_2 ),
       .io_outPort_1( Switch_34_io_outPort_1 ),
       .io_outPort_0( Switch_34_io_outPort_0 ),
       .io_deqValid( Switch_34_io_deqValid ),
       .io_enqRdy( Switch_34_io_enqRdy ),
       .io_deqRdy( T31 ),
       .io_enqValid( T21 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( Switch_35_io_enqOR ),
       .io_enqOR( Switch_34_io_enqOR ),
       .io_deqRdyOut( T18 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_34.io_inPort_7 = {2{$random}};
    assign Switch_34.io_inPort_4 = {2{$random}};
// synthesis translate_on
`endif
  Switch_5 Switch_35(.clk(clk), .reset(reset),
       //.io_inPort_7(  )
       .io_inPort_6( CU_24_io_out ),
       //.io_inPort_5(  )
       //.io_inPort_4(  )
       .io_inPort_3( Switch_34_io_outPort_1 ),
       .io_inPort_2( Switch_29_io_outPort_0 ),
       .io_inPort_1( io_inData_10 ),
       //.io_inPort_0(  )
       //.io_outPort_7(  )
       .io_outPort_6( Switch_35_io_outPort_6 ),
       //.io_outPort_5(  )
       //.io_outPort_4(  )
       .io_outPort_3( Switch_35_io_outPort_3 ),
       .io_outPort_2( Switch_35_io_outPort_2 ),
       .io_outPort_1( Switch_35_io_outPort_1 ),
       //.io_outPort_0(  )
       .io_deqValid( Switch_35_io_deqValid ),
       .io_enqRdy( Switch_35_io_enqRdy ),
       .io_deqRdy( T10 ),
       .io_enqValid( T2 ),
       //.io_outConfigData(  )
       //.io_outCUConfig(  )
       .io_deqOR( 1'h0 ),
       .io_enqOR( Switch_35_io_enqOR ),
       .io_deqRdyOut( T0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Switch_35.io_inPort_7 = {2{$random}};
    assign Switch_35.io_inPort_5 = {2{$random}};
    assign Switch_35.io_inPort_4 = {2{$random}};
    assign Switch_35.io_inPort_0 = {2{$random}};
// synthesis translate_on
`endif
endmodule

