module controllerConfigure_0(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_outConfig,
    output io_outValid,
    output io_computeCtrl,
    output io_computeCtrlValid
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  reg [31:0] inDataReg;
  wire[31:0] T30;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inDataReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_computeCtrlValid = T0;
  assign T0 = T21 ? 1'h0 : T1;
  assign T1 = T18 ? 1'h1 : T2;
  assign T2 = T13 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : 1'h0;
  assign T4 = T11 & T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 2'h0;
  assign T7 = inDataReg[5'h1f:5'h1e];
  assign T30 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inDataReg;
  assign T9 = T10 == 1'h1;
  assign T10 = inDataReg[1'h0:1'h0];
  assign T11 = T12 == 1'h0;
  assign T12 = inDataReg[5'h1f:5'h1f];
  assign T13 = T11 & T14;
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h102;
  assign T16 = inDataReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T11 & T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T5 | T15;
  assign T21 = T11 ^ 1'h1;
  assign io_computeCtrl = T22;
  assign T22 = T21 ? 1'h0 : T23;
  assign T23 = T18 ? 1'h0 : T24;
  assign T24 = T13 ? 1'h0 : T25;
  assign T25 = T4 ? 1'h1 : 1'h0;
  assign io_outValid = T26;
  assign T26 = T21 ? 1'h0 : T27;
  assign T27 = T18 ? 1'h0 : T28;
  assign T28 = T13 ? 1'h1 : T29;
  assign T29 = T4 ? 1'h0 : 1'h0;
  assign io_outConfig = inDataReg;

  always @(posedge clk) begin
    if(reset) begin
      inDataReg <= 32'h0;
    end else if(io_inValid) begin
      inDataReg <= io_inConfig;
    end
  end
endmodule

module fabInSeqCtrl(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[8:0] io_seqMemAddr,
    output io_seqMemAddrValid,
    input  io_seqProceed,
    output io_computeDone
);

  wire T0;
  reg  computeEnable;
  wire T119;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[514:0] lastAddr;
  wire[514:0] T120;
  wire[513:0] T7;
  wire[513:0] T121;
  reg [8:0] epilogueDepth;
  wire[8:0] T122;
  wire[8:0] T8;
  wire[8:0] T123;
  wire[6:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire[9:0] T22;
  wire[513:0] ssEnd;
  wire[513:0] T124;
  wire[8:0] T23;
  reg [8:0] steadyStateDepth;
  wire[8:0] T125;
  wire[9:0] T126;
  wire[9:0] T24;
  wire[9:0] T127;
  wire[9:0] T25;
  wire T26;
  reg [8:0] prologueDepth;
  wire[8:0] T128;
  wire[8:0] T27;
  wire[8:0] T129;
  wire[6:0] T28;
  wire startComputeValid;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire computeDone;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[514:0] T37;
  wire[514:0] T130;
  reg [511:0] seqMemAddr;
  wire[511:0] T131;
  wire[513:0] T132;
  wire[513:0] T38;
  wire[513:0] T39;
  wire[513:0] T133;
  wire[511:0] T40;
  wire[511:0] T41;
  wire[511:0] T42;
  wire T43;
  wire T44;
  wire nextRequest;
  wire T45;
  wire T46;
  wire T47;
  wire[511:0] T134;
  wire T48;
  wire T49;
  wire T50;
  reg [8:0] epilogueSpill;
  wire[8:0] T135;
  wire[9:0] T136;
  wire[9:0] T51;
  wire[9:0] T137;
  wire[9:0] T52;
  wire T53;
  wire[31:0] T54;
  reg [31:0] iterCount;
  wire[31:0] T138;
  wire[31:0] T55;
  wire[31:0] T139;
  wire[18:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire[2:0] T60;
  wire T61;
  reg [31:0] currentIter;
  wire[31:0] T140;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire T65;
  wire T66;
  wire[513:0] T67;
  wire[513:0] T141;
  wire T68;
  wire T69;
  wire[511:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[513:0] T77;
  wire[513:0] T142;
  wire T78;
  wire T79;
  wire[513:0] T143;
  wire[511:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[31:0] T91;
  wire T92;
  wire[514:0] T93;
  wire[514:0] T144;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[513:0] T101;
  wire[513:0] spillEndAddr;
  wire[513:0] T145;
  wire[8:0] T102;
  wire[513:0] T146;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire resetComputeValid;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[8:0] T147;
  wire[511:0] T117;
  wire[511:0] T118;
  wire fabInSeqCtrlConfigure_io_computeCtrl;
  wire fabInSeqCtrlConfigure_io_computeCtrlValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    computeEnable = {1{$random}};
    epilogueDepth = {1{$random}};
    steadyStateDepth = {1{$random}};
    prologueDepth = {1{$random}};
    seqMemAddr = {16{$random}};
    epilogueSpill = {1{$random}};
    iterCount = {1{$random}};
    currentIter = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_computeDone = T0;
  assign T0 = computeEnable ^ 1'h1;
  assign T119 = reset ? 1'h0 : T1;
  assign T1 = T113 ? 1'h0 : T2;
  assign T2 = T110 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : computeEnable;
  assign T4 = T32 & T5;
  assign T5 = startComputeValid & T6;
  assign T6 = lastAddr != 515'h0;
  assign lastAddr = T120;
  assign T120 = {1'h0, T7};
  assign T7 = ssEnd + T121;
  assign T121 = {505'h0, epilogueDepth};
  assign T122 = reset ? 9'h0 : T8;
  assign T8 = T10 ? T123 : epilogueDepth;
  assign T123 = {2'h0, T9};
  assign T9 = io_inConfig[3'h6:1'h0];
  assign T10 = T17 & T11;
  assign T11 = T14 & T12;
  assign T12 = T13 == 1'h1;
  assign T13 = io_inConfig[5'h11:5'h11];
  assign T14 = T15 ^ 1'h1;
  assign T15 = T16 == 1'h0;
  assign T16 = io_inConfig[5'h11:5'h11];
  assign T17 = T20 & T18;
  assign T18 = T19 == 3'h0;
  assign T19 = io_inConfig[5'h15:5'h13];
  assign T20 = io_inValid & T21;
  assign T21 = T22 == 10'h103;
  assign T22 = io_inConfig[5'h1f:5'h16];
  assign ssEnd = T124;
  assign T124 = {505'h0, T23};
  assign T23 = prologueDepth + steadyStateDepth;
  assign T125 = T126[4'h8:1'h0];
  assign T126 = reset ? 10'h0 : T24;
  assign T24 = T26 ? T25 : T127;
  assign T127 = {1'h0, steadyStateDepth};
  assign T25 = io_inConfig[5'h10:3'h7];
  assign T26 = T17 & T15;
  assign T128 = reset ? 9'h0 : T27;
  assign T27 = T26 ? T129 : prologueDepth;
  assign T129 = {2'h0, T28};
  assign T28 = io_inConfig[3'h6:1'h0];
  assign startComputeValid = T29;
  assign T29 = T31 ? 1'h0 : T30;
  assign T30 = fabInSeqCtrlConfigure_io_computeCtrlValid & fabInSeqCtrlConfigure_io_computeCtrl;
  assign T31 = fabInSeqCtrlConfigure_io_computeCtrlValid ^ 1'h1;
  assign T32 = T106 | computeDone;
  assign computeDone = T33;
  assign T33 = T103 ? T98 : T34;
  assign T34 = T94 ? T89 : T35;
  assign T35 = T84 ? T36 : 1'h0;
  assign T36 = T130 == T37;
  assign T37 = lastAddr - 515'h1;
  assign T130 = {3'h0, seqMemAddr};
  assign T131 = T132[9'h1ff:1'h0];
  assign T132 = reset ? 514'h0 : T38;
  assign T38 = T81 ? T143 : T39;
  assign T39 = T73 ? ssEnd : T133;
  assign T133 = {2'h0, T40};
  assign T40 = T71 ? T70 : T41;
  assign T41 = T48 ? T134 : T42;
  assign T42 = T43 ? 512'h0 : seqMemAddr;
  assign T43 = T44 & startComputeValid;
  assign T44 = startComputeValid | nextRequest;
  assign nextRequest = T45;
  assign T45 = T47 ? 1'h0 : T46;
  assign T46 = io_seqProceed & computeEnable;
  assign T47 = T46 ^ 1'h1;
  assign T134 = {503'h0, prologueDepth};
  assign T48 = T65 & T49;
  assign T49 = T53 | T50;
  assign T50 = epilogueSpill != 9'h0;
  assign T135 = T136[4'h8:1'h0];
  assign T136 = reset ? 10'h0 : T51;
  assign T51 = T10 ? T52 : T137;
  assign T137 = {1'h0, epilogueSpill};
  assign T52 = io_inConfig[5'h10:3'h7];
  assign T53 = currentIter < T54;
  assign T54 = iterCount - 32'h1;
  assign T138 = reset ? 32'h0 : T55;
  assign T55 = T57 ? T139 : iterCount;
  assign T139 = {13'h0, T56};
  assign T56 = io_inConfig[5'h12:1'h0];
  assign T57 = T20 & T58;
  assign T58 = T61 & T59;
  assign T59 = T60 == 3'h1;
  assign T60 = io_inConfig[5'h15:5'h13];
  assign T61 = T18 ^ 1'h1;
  assign T140 = reset ? 32'h0 : T62;
  assign T62 = T48 ? T64 : T63;
  assign T63 = T43 ? 32'h0 : currentIter;
  assign T64 = currentIter + 32'h1;
  assign T65 = T68 & T66;
  assign T66 = T141 == T67;
  assign T67 = ssEnd - 514'h1;
  assign T141 = {2'h0, seqMemAddr};
  assign T68 = T44 & T69;
  assign T69 = startComputeValid ^ 1'h1;
  assign T70 = seqMemAddr + 512'h1;
  assign T71 = T65 & T72;
  assign T72 = T49 ^ 1'h1;
  assign T73 = T68 & T74;
  assign T74 = T79 & T75;
  assign T75 = T78 & T76;
  assign T76 = T142 == T77;
  assign T77 = ssEnd - 514'h1;
  assign T142 = {2'h0, seqMemAddr};
  assign T78 = currentIter == iterCount;
  assign T79 = T66 ^ 1'h1;
  assign T143 = {2'h0, T80};
  assign T80 = seqMemAddr + 512'h1;
  assign T81 = T68 & T82;
  assign T82 = T83 ^ 1'h1;
  assign T83 = T66 | T75;
  assign T84 = T88 & T85;
  assign T85 = T87 & T86;
  assign T86 = steadyStateDepth == 9'h0;
  assign T87 = epilogueDepth != 9'h0;
  assign T88 = computeEnable & nextRequest;
  assign T89 = T92 & T90;
  assign T90 = T91 == iterCount;
  assign T91 = currentIter + 32'h1;
  assign T92 = T144 == T93;
  assign T93 = lastAddr - 515'h1;
  assign T144 = {3'h0, seqMemAddr};
  assign T94 = T88 & T95;
  assign T95 = T97 & T96;
  assign T96 = epilogueSpill == 9'h0;
  assign T97 = T85 ^ 1'h1;
  assign T98 = T100 & T99;
  assign T99 = currentIter == iterCount;
  assign T100 = T146 == T101;
  assign T101 = spillEndAddr - 514'h1;
  assign spillEndAddr = T145;
  assign T145 = {505'h0, T102};
  assign T102 = prologueDepth + epilogueSpill;
  assign T146 = {2'h0, seqMemAddr};
  assign T103 = T88 & T104;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T85 | T96;
  assign T106 = startComputeValid | resetComputeValid;
  assign resetComputeValid = T107;
  assign T107 = T31 ? 1'h0 : T108;
  assign T108 = fabInSeqCtrlConfigure_io_computeCtrlValid & T109;
  assign T109 = fabInSeqCtrlConfigure_io_computeCtrl ^ 1'h1;
  assign T110 = T32 & T111;
  assign T111 = T112 & resetComputeValid;
  assign T112 = T5 ^ 1'h1;
  assign T113 = T32 & T114;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T5 | resetComputeValid;
  assign io_seqMemAddrValid = T116;
  assign T116 = T46 ? 1'h1 : 1'h0;
  assign io_seqMemAddr = T147;
  assign T147 = T117[4'h8:1'h0];
  assign T117 = T46 ? seqMemAddr : T118;
  assign T118 = T44 ? seqMemAddr : seqMemAddr;
  controllerConfigure_0 fabInSeqCtrlConfigure(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       //.io_outConfig(  )
       //.io_outValid(  )
       .io_computeCtrl( fabInSeqCtrlConfigure_io_computeCtrl ),
       .io_computeCtrlValid( fabInSeqCtrlConfigure_io_computeCtrlValid )
  );

  always @(posedge clk) begin
    if(reset) begin
      computeEnable <= 1'h0;
    end else if(T113) begin
      computeEnable <= 1'h0;
    end else if(T110) begin
      computeEnable <= 1'h0;
    end else if(T4) begin
      computeEnable <= 1'h1;
    end
    if(reset) begin
      epilogueDepth <= 9'h0;
    end else if(T10) begin
      epilogueDepth <= T123;
    end
    steadyStateDepth <= T125;
    if(reset) begin
      prologueDepth <= 9'h0;
    end else if(T26) begin
      prologueDepth <= T129;
    end
    seqMemAddr <= T131;
    epilogueSpill <= T135;
    if(reset) begin
      iterCount <= 32'h0;
    end else if(T57) begin
      iterCount <= T139;
    end
    if(reset) begin
      currentIter <= 32'h0;
    end else if(T48) begin
      currentIter <= T64;
    end else if(T43) begin
      currentIter <= 32'h0;
    end
  end
endmodule

module customReg_0(input clk,
    input [88:0] io_inData,
    output[88:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [8:0] io_readAddr,
    input [8:0] io_writeAddr
);

  wire[88:0] T0;
  reg [88:0] ram [511:0];
  wire[88:0] T1;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 512; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];

  always @(posedge clk) begin
    if (io_writeEn)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module fifo_6(input clk, input reset,
    input [43:0] io_enqData,
    output[43:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg  deqPtr;
  wire T21;
  wire T2;
  wire T3;
  wire deqPtrInc;
  wire T4;
  wire doDeq;
  wire T5;
  reg  enqPtr;
  wire T22;
  wire T6;
  wire T7;
  wire enqPtrInc;
  wire T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[43:0] T19;
  reg [43:0] fifoMem [1:0];
  wire[43:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = io_rst ? 1'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 2'h2;
  assign T4 = deqPtr + 1'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 1'h0 : T6;
  assign T6 = io_rst ? 1'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 2'h2;
  assign T8 = enqPtr + 1'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(io_rst) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(io_rst) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module customReg_5(input clk,
    input [31:0] io_inData,
    output[31:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [5:0] io_readAddr,
    input [5:0] io_writeAddr
);

  wire[31:0] T0;
  reg [31:0] ram [63:0];
  wire[31:0] T1;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 64; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];

  always @(posedge clk) begin
    if (io_writeEn)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module memoryBank(input clk, input reset,
    input [31:0] io_inData,
    output[31:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    output io_writeSuccess,
    output io_readSuccess,
    input  io_doInvalidate,
    output io_isValid,
    output io_isWriteLoadRdy,
    output io_isWriteFabricRdy,
    input [5:0] io_readAddr,
    input [5:0] io_writeAddr,
    input [5:0] io_writeLoadAddr,
    input [5:0] io_writeFabricAddr,
    input  io_rst
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[5:0] T5;
  wire[5:0] T6;
  wire T7;
  reg [63:0] validBit;
  wire[63:0] T76;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T11;
  wire[63:0] T12;
  wire[63:0] T13;
  wire[63:0] T14;
  wire[63:0] T15;
  wire[63:0] T77;
  wire T16;
  wire T17;
  wire[63:0] T18;
  wire[63:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[5:0] T25;
  wire[5:0] T26;
  wire T27;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] T78;
  wire T33;
  wire T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[5:0] T46;
  wire[5:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[5:0] T58;
  wire[5:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[5:0] T70;
  wire[5:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[31:0] memoryClass_io_outData;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    validBit = {2{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_writeEn & T1;
  assign T1 = ~ T2;
  assign T2 = T7 & T3;
  assign T3 = T4 - 1'h1;
  assign T4 = 1'h1 << T5;
  assign T5 = T6 + 6'h1;
  assign T6 = io_writeAddr - io_writeAddr;
  assign T7 = validBit >> io_writeAddr;
  assign T76 = reset ? 64'h0 : T8;
  assign T8 = T37 ? T28 : T9;
  assign T9 = T20 ? T11 : T10;
  assign T10 = io_rst ? 64'h0 : validBit;
  assign T11 = T18 | T12;
  assign T12 = T77 & T13;
  assign T13 = T15 | T14;
  assign T14 = validBit ^ validBit;
  assign T15 = 1'h1 << io_readAddr;
  assign T77 = T16 ? 64'hffffffffffffffff : 64'h0;
  assign T16 = T17;
  assign T17 = 1'h0;
  assign T18 = T10 & T19;
  assign T19 = ~ T13;
  assign T20 = T21 & io_doInvalidate;
  assign T21 = io_readEn & T22;
  assign T22 = T27 & T23;
  assign T23 = T24 - 1'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = T26 + 6'h1;
  assign T26 = io_readAddr - io_readAddr;
  assign T27 = validBit >> io_readAddr;
  assign T28 = T35 | T29;
  assign T29 = T78 & T30;
  assign T30 = T32 | T31;
  assign T31 = validBit ^ validBit;
  assign T32 = 1'h1 << io_writeAddr;
  assign T78 = T33 ? 64'hffffffffffffffff : 64'h0;
  assign T33 = T34;
  assign T34 = 1'h1;
  assign T35 = T9 & T36;
  assign T36 = ~ T30;
  assign T37 = T41 | T38;
  assign T38 = T39 & io_doInvalidate;
  assign T39 = T40 & io_readEn;
  assign T40 = io_readAddr == io_writeAddr;
  assign T41 = io_writeEn & T42;
  assign T42 = ~ T43;
  assign T43 = T48 & T44;
  assign T44 = T45 - 1'h1;
  assign T45 = 1'h1 << T46;
  assign T46 = T47 + 6'h1;
  assign T47 = io_writeAddr - io_writeAddr;
  assign T48 = validBit >> io_writeAddr;
  assign io_isWriteFabricRdy = T49;
  assign T49 = T50 ? 1'h1 : 1'h0;
  assign T50 = T54 | T51;
  assign T51 = T52 & io_doInvalidate;
  assign T52 = T53 & io_readEn;
  assign T53 = io_readAddr == io_writeFabricAddr;
  assign T54 = ~ T55;
  assign T55 = T60 & T56;
  assign T56 = T57 - 1'h1;
  assign T57 = 1'h1 << T58;
  assign T58 = T59 + 6'h1;
  assign T59 = io_writeFabricAddr - io_writeFabricAddr;
  assign T60 = validBit >> io_writeFabricAddr;
  assign io_isWriteLoadRdy = T61;
  assign T61 = T62 ? 1'h1 : 1'h0;
  assign T62 = T66 | T63;
  assign T63 = T64 & io_doInvalidate;
  assign T64 = T65 & io_readEn;
  assign T65 = io_readAddr == io_writeLoadAddr;
  assign T66 = ~ T67;
  assign T67 = T72 & T68;
  assign T68 = T69 - 1'h1;
  assign T69 = 1'h1 << T70;
  assign T70 = T71 + 6'h1;
  assign T71 = io_writeLoadAddr - io_writeLoadAddr;
  assign T72 = validBit >> io_writeLoadAddr;
  assign io_isValid = T73;
  assign T73 = T21 ? 1'h1 : 1'h0;
  assign io_readSuccess = T74;
  assign T74 = T21 ? 1'h1 : 1'h0;
  assign io_writeSuccess = T75;
  assign T75 = T37 ? 1'h1 : 1'h0;
  assign io_outData = memoryClass_io_outData;
  customReg_5 memoryClass(.clk(clk),
       .io_inData( io_inData ),
       .io_outData( memoryClass_io_outData ),
       .io_readEn( io_readEn ),
       .io_writeEn( T0 ),
       .io_readAddr( io_readAddr ),
       .io_writeAddr( io_writeAddr )
  );

  always @(posedge clk) begin
    if(reset) begin
      validBit <= 64'h0;
    end else if(T37) begin
      validBit <= T28;
    end else if(T20) begin
      validBit <= T11;
    end else if(io_rst) begin
      validBit <= 64'h0;
    end
  end
endmodule

module controllerLocalStorage(input clk, input reset,
    input [37:0] io_inDataLoad_7,
    input [37:0] io_inDataLoad_6,
    input [37:0] io_inDataLoad_5,
    input [37:0] io_inDataLoad_4,
    input [37:0] io_inDataLoad_3,
    input [37:0] io_inDataLoad_2,
    input [37:0] io_inDataLoad_1,
    input [37:0] io_inDataLoad_0,
    input [37:0] io_inDataFabric_7,
    input [37:0] io_inDataFabric_6,
    input [37:0] io_inDataFabric_5,
    input [37:0] io_inDataFabric_4,
    input [37:0] io_inDataFabric_3,
    input [37:0] io_inDataFabric_2,
    input [37:0] io_inDataFabric_1,
    input [37:0] io_inDataFabric_0,
    output[37:0] io_outData_7,
    output[37:0] io_outData_6,
    output[37:0] io_outData_5,
    output[37:0] io_outData_4,
    output[37:0] io_outData_3,
    output[37:0] io_outData_2,
    output[37:0] io_outData_1,
    output[37:0] io_outData_0,
    output io_isReadValid_7,
    output io_isReadValid_6,
    output io_isReadValid_5,
    output io_isReadValid_4,
    output io_isReadValid_3,
    output io_isReadValid_2,
    output io_isReadValid_1,
    output io_isReadValid_0,
    input [5:0] io_readAddr_7,
    input [5:0] io_readAddr_6,
    input [5:0] io_readAddr_5,
    input [5:0] io_readAddr_4,
    input [5:0] io_readAddr_3,
    input [5:0] io_readAddr_2,
    input [5:0] io_readAddr_1,
    input [5:0] io_readAddr_0,
    input  io_readEn_7,
    input  io_readEn_6,
    input  io_readEn_5,
    input  io_readEn_4,
    input  io_readEn_3,
    input  io_readEn_2,
    input  io_readEn_1,
    input  io_readEn_0,
    input  io_doInvalidate_7,
    input  io_doInvalidate_6,
    input  io_doInvalidate_5,
    input  io_doInvalidate_4,
    input  io_doInvalidate_3,
    input  io_doInvalidate_2,
    input  io_doInvalidate_1,
    input  io_doInvalidate_0,
    output io_readSuccess_7,
    output io_readSuccess_6,
    output io_readSuccess_5,
    output io_readSuccess_4,
    output io_readSuccess_3,
    output io_readSuccess_2,
    output io_readSuccess_1,
    output io_readSuccess_0,
    output io_writeSuccess_7,
    output io_writeSuccess_6,
    output io_writeSuccess_5,
    output io_writeSuccess_4,
    output io_writeSuccess_3,
    output io_writeSuccess_2,
    output io_writeSuccess_1,
    output io_writeSuccess_0,
    output io_enqRdyLoad_7,
    output io_enqRdyLoad_6,
    output io_enqRdyLoad_5,
    output io_enqRdyLoad_4,
    output io_enqRdyLoad_3,
    output io_enqRdyLoad_2,
    output io_enqRdyLoad_1,
    output io_enqRdyLoad_0,
    output io_enqRdyFabric_7,
    output io_enqRdyFabric_6,
    output io_enqRdyFabric_5,
    output io_enqRdyFabric_4,
    output io_enqRdyFabric_3,
    output io_enqRdyFabric_2,
    output io_enqRdyFabric_1,
    output io_enqRdyFabric_0,
    input  io_enqValidLoad_7,
    input  io_enqValidLoad_6,
    input  io_enqValidLoad_5,
    input  io_enqValidLoad_4,
    input  io_enqValidLoad_3,
    input  io_enqValidLoad_2,
    input  io_enqValidLoad_1,
    input  io_enqValidLoad_0,
    input  io_enqValidFabric_7,
    input  io_enqValidFabric_6,
    input  io_enqValidFabric_5,
    input  io_enqValidFabric_4,
    input  io_enqValidFabric_3,
    input  io_enqValidFabric_2,
    input  io_enqValidFabric_1,
    input  io_enqValidFabric_0,
    input  io_rst
);

  wire[5:0] T0;
  wire[5:0] T1;
  wire[5:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire[5:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire[31:0] T176;
  wire[37:0] T14;
  wire[37:0] T15;
  wire[37:0] T16;
  wire[37:0] T17;
  wire[5:0] T18;
  wire[5:0] T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire[5:0] T22;
  wire T23;
  wire T24;
  wire[5:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[31:0] T177;
  wire[37:0] T32;
  wire[37:0] T33;
  wire[37:0] T34;
  wire[37:0] T35;
  wire[5:0] T36;
  wire[5:0] T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire T41;
  wire T42;
  wire[5:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[31:0] T178;
  wire[37:0] T50;
  wire[37:0] T51;
  wire[37:0] T52;
  wire[37:0] T53;
  wire[5:0] T54;
  wire[5:0] T55;
  wire[5:0] T56;
  wire[5:0] T57;
  wire[5:0] T58;
  wire T59;
  wire T60;
  wire[5:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[31:0] T179;
  wire[37:0] T68;
  wire[37:0] T69;
  wire[37:0] T70;
  wire[37:0] T71;
  wire[5:0] T72;
  wire[5:0] T73;
  wire[5:0] T74;
  wire[5:0] T75;
  wire[5:0] T76;
  wire T77;
  wire T78;
  wire[5:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[31:0] T180;
  wire[37:0] T86;
  wire[37:0] T87;
  wire[37:0] T88;
  wire[37:0] T89;
  wire[5:0] T90;
  wire[5:0] T91;
  wire[5:0] T92;
  wire[5:0] T93;
  wire[5:0] T94;
  wire T95;
  wire T96;
  wire[5:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[31:0] T181;
  wire[37:0] T104;
  wire[37:0] T105;
  wire[37:0] T106;
  wire[37:0] T107;
  wire[5:0] T108;
  wire[5:0] T109;
  wire[5:0] T110;
  wire[5:0] T111;
  wire[5:0] T112;
  wire T113;
  wire T114;
  wire[5:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[31:0] T182;
  wire[37:0] T122;
  wire[37:0] T123;
  wire[37:0] T124;
  wire[37:0] T125;
  wire[5:0] T126;
  wire[5:0] T127;
  wire[5:0] T128;
  wire[5:0] T129;
  wire[5:0] T130;
  wire T131;
  wire T132;
  wire[5:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[31:0] T183;
  wire[37:0] T140;
  wire[37:0] T141;
  wire[37:0] T142;
  wire[37:0] T143;
  wire T144;
  wire[43:0] T184;
  wire T145;
  wire[43:0] T185;
  wire T146;
  wire[43:0] T186;
  wire T147;
  wire[43:0] T187;
  wire T148;
  wire[43:0] T188;
  wire T149;
  wire[43:0] T189;
  wire T150;
  wire[43:0] T190;
  wire T151;
  wire[43:0] T191;
  wire T152;
  wire[43:0] T192;
  wire T153;
  wire[43:0] T193;
  wire T154;
  wire[43:0] T194;
  wire T155;
  wire[43:0] T195;
  wire T156;
  wire[43:0] T196;
  wire T157;
  wire[43:0] T197;
  wire T158;
  wire[43:0] T198;
  wire T159;
  wire[43:0] T199;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[37:0] T200;
  wire[37:0] T201;
  wire[37:0] T202;
  wire[37:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[37:0] T206;
  wire[37:0] T207;
  wire[43:0] fifo_io_deqData;
  wire fifo_io_enqRdy;
  wire fifo_io_deqValid;
  wire[43:0] fifo_1_io_deqData;
  wire fifo_1_io_enqRdy;
  wire fifo_1_io_deqValid;
  wire[43:0] fifo_2_io_deqData;
  wire fifo_2_io_enqRdy;
  wire fifo_2_io_deqValid;
  wire[43:0] fifo_3_io_deqData;
  wire fifo_3_io_enqRdy;
  wire fifo_3_io_deqValid;
  wire[43:0] fifo_4_io_deqData;
  wire fifo_4_io_enqRdy;
  wire fifo_4_io_deqValid;
  wire[43:0] fifo_5_io_deqData;
  wire fifo_5_io_enqRdy;
  wire fifo_5_io_deqValid;
  wire[43:0] fifo_6_io_deqData;
  wire fifo_6_io_enqRdy;
  wire fifo_6_io_deqValid;
  wire[43:0] fifo_7_io_deqData;
  wire fifo_7_io_enqRdy;
  wire fifo_7_io_deqValid;
  wire[43:0] fifo_8_io_deqData;
  wire fifo_8_io_enqRdy;
  wire fifo_8_io_deqValid;
  wire[43:0] fifo_9_io_deqData;
  wire fifo_9_io_enqRdy;
  wire fifo_9_io_deqValid;
  wire[43:0] fifo_10_io_deqData;
  wire fifo_10_io_enqRdy;
  wire fifo_10_io_deqValid;
  wire[43:0] fifo_11_io_deqData;
  wire fifo_11_io_enqRdy;
  wire fifo_11_io_deqValid;
  wire[43:0] fifo_12_io_deqData;
  wire fifo_12_io_enqRdy;
  wire fifo_12_io_deqValid;
  wire[43:0] fifo_13_io_deqData;
  wire fifo_13_io_enqRdy;
  wire fifo_13_io_deqValid;
  wire[43:0] fifo_14_io_deqData;
  wire fifo_14_io_enqRdy;
  wire fifo_14_io_deqValid;
  wire[43:0] fifo_15_io_deqData;
  wire fifo_15_io_enqRdy;
  wire fifo_15_io_deqValid;
  wire[31:0] memoryBank_io_outData;
  wire memoryBank_io_writeSuccess;
  wire memoryBank_io_readSuccess;
  wire memoryBank_io_isValid;
  wire memoryBank_io_isWriteLoadRdy;
  wire memoryBank_io_isWriteFabricRdy;
  wire[31:0] memoryBank_1_io_outData;
  wire memoryBank_1_io_writeSuccess;
  wire memoryBank_1_io_readSuccess;
  wire memoryBank_1_io_isValid;
  wire memoryBank_1_io_isWriteLoadRdy;
  wire memoryBank_1_io_isWriteFabricRdy;
  wire[31:0] memoryBank_2_io_outData;
  wire memoryBank_2_io_writeSuccess;
  wire memoryBank_2_io_readSuccess;
  wire memoryBank_2_io_isValid;
  wire memoryBank_2_io_isWriteLoadRdy;
  wire memoryBank_2_io_isWriteFabricRdy;
  wire[31:0] memoryBank_3_io_outData;
  wire memoryBank_3_io_writeSuccess;
  wire memoryBank_3_io_readSuccess;
  wire memoryBank_3_io_isValid;
  wire memoryBank_3_io_isWriteLoadRdy;
  wire memoryBank_3_io_isWriteFabricRdy;
  wire[31:0] memoryBank_4_io_outData;
  wire memoryBank_4_io_writeSuccess;
  wire memoryBank_4_io_readSuccess;
  wire memoryBank_4_io_isValid;
  wire memoryBank_4_io_isWriteLoadRdy;
  wire memoryBank_4_io_isWriteFabricRdy;
  wire[31:0] memoryBank_5_io_outData;
  wire memoryBank_5_io_writeSuccess;
  wire memoryBank_5_io_readSuccess;
  wire memoryBank_5_io_isValid;
  wire memoryBank_5_io_isWriteLoadRdy;
  wire memoryBank_5_io_isWriteFabricRdy;
  wire[31:0] memoryBank_6_io_outData;
  wire memoryBank_6_io_writeSuccess;
  wire memoryBank_6_io_readSuccess;
  wire memoryBank_6_io_isValid;
  wire memoryBank_6_io_isWriteLoadRdy;
  wire memoryBank_6_io_isWriteFabricRdy;
  wire[31:0] memoryBank_7_io_outData;
  wire memoryBank_7_io_writeSuccess;
  wire memoryBank_7_io_readSuccess;
  wire memoryBank_7_io_isValid;
  wire memoryBank_7_io_isWriteLoadRdy;
  wire memoryBank_7_io_isWriteFabricRdy;


  assign T0 = fifo_15_io_deqData[6'h2b:6'h26];
  assign T1 = fifo_7_io_deqData[6'h2b:6'h26];
  assign T2 = T8 ? T7 : T3;
  assign T3 = T5 ? T4 : 6'h0;
  assign T4 = fifo_7_io_deqData[6'h2b:6'h26];
  assign T5 = T6 & memoryBank_7_io_isWriteLoadRdy;
  assign T6 = fifo_7_io_deqValid;
  assign T7 = fifo_15_io_deqData[6'h2b:6'h26];
  assign T8 = T11 & T9;
  assign T9 = T10 & memoryBank_7_io_isWriteFabricRdy;
  assign T10 = fifo_15_io_deqValid;
  assign T11 = T5 ^ 1'h1;
  assign T12 = T8 ? 1'h1 : T13;
  assign T13 = T5 ? 1'h1 : 1'h0;
  assign T176 = T14[5'h1f:1'h0];
  assign T14 = T8 ? T17 : T15;
  assign T15 = T5 ? T16 : 38'h0;
  assign T16 = fifo_7_io_deqData[6'h25:1'h0];
  assign T17 = fifo_15_io_deqData[6'h25:1'h0];
  assign T18 = fifo_14_io_deqData[6'h2b:6'h26];
  assign T19 = fifo_6_io_deqData[6'h2b:6'h26];
  assign T20 = T26 ? T25 : T21;
  assign T21 = T23 ? T22 : 6'h0;
  assign T22 = fifo_6_io_deqData[6'h2b:6'h26];
  assign T23 = T24 & memoryBank_6_io_isWriteLoadRdy;
  assign T24 = fifo_6_io_deqValid;
  assign T25 = fifo_14_io_deqData[6'h2b:6'h26];
  assign T26 = T29 & T27;
  assign T27 = T28 & memoryBank_6_io_isWriteFabricRdy;
  assign T28 = fifo_14_io_deqValid;
  assign T29 = T23 ^ 1'h1;
  assign T30 = T26 ? 1'h1 : T31;
  assign T31 = T23 ? 1'h1 : 1'h0;
  assign T177 = T32[5'h1f:1'h0];
  assign T32 = T26 ? T35 : T33;
  assign T33 = T23 ? T34 : 38'h0;
  assign T34 = fifo_6_io_deqData[6'h25:1'h0];
  assign T35 = fifo_14_io_deqData[6'h25:1'h0];
  assign T36 = fifo_13_io_deqData[6'h2b:6'h26];
  assign T37 = fifo_5_io_deqData[6'h2b:6'h26];
  assign T38 = T44 ? T43 : T39;
  assign T39 = T41 ? T40 : 6'h0;
  assign T40 = fifo_5_io_deqData[6'h2b:6'h26];
  assign T41 = T42 & memoryBank_5_io_isWriteLoadRdy;
  assign T42 = fifo_5_io_deqValid;
  assign T43 = fifo_13_io_deqData[6'h2b:6'h26];
  assign T44 = T47 & T45;
  assign T45 = T46 & memoryBank_5_io_isWriteFabricRdy;
  assign T46 = fifo_13_io_deqValid;
  assign T47 = T41 ^ 1'h1;
  assign T48 = T44 ? 1'h1 : T49;
  assign T49 = T41 ? 1'h1 : 1'h0;
  assign T178 = T50[5'h1f:1'h0];
  assign T50 = T44 ? T53 : T51;
  assign T51 = T41 ? T52 : 38'h0;
  assign T52 = fifo_5_io_deqData[6'h25:1'h0];
  assign T53 = fifo_13_io_deqData[6'h25:1'h0];
  assign T54 = fifo_12_io_deqData[6'h2b:6'h26];
  assign T55 = fifo_4_io_deqData[6'h2b:6'h26];
  assign T56 = T62 ? T61 : T57;
  assign T57 = T59 ? T58 : 6'h0;
  assign T58 = fifo_4_io_deqData[6'h2b:6'h26];
  assign T59 = T60 & memoryBank_4_io_isWriteLoadRdy;
  assign T60 = fifo_4_io_deqValid;
  assign T61 = fifo_12_io_deqData[6'h2b:6'h26];
  assign T62 = T65 & T63;
  assign T63 = T64 & memoryBank_4_io_isWriteFabricRdy;
  assign T64 = fifo_12_io_deqValid;
  assign T65 = T59 ^ 1'h1;
  assign T66 = T62 ? 1'h1 : T67;
  assign T67 = T59 ? 1'h1 : 1'h0;
  assign T179 = T68[5'h1f:1'h0];
  assign T68 = T62 ? T71 : T69;
  assign T69 = T59 ? T70 : 38'h0;
  assign T70 = fifo_4_io_deqData[6'h25:1'h0];
  assign T71 = fifo_12_io_deqData[6'h25:1'h0];
  assign T72 = fifo_11_io_deqData[6'h2b:6'h26];
  assign T73 = fifo_3_io_deqData[6'h2b:6'h26];
  assign T74 = T80 ? T79 : T75;
  assign T75 = T77 ? T76 : 6'h0;
  assign T76 = fifo_3_io_deqData[6'h2b:6'h26];
  assign T77 = T78 & memoryBank_3_io_isWriteLoadRdy;
  assign T78 = fifo_3_io_deqValid;
  assign T79 = fifo_11_io_deqData[6'h2b:6'h26];
  assign T80 = T83 & T81;
  assign T81 = T82 & memoryBank_3_io_isWriteFabricRdy;
  assign T82 = fifo_11_io_deqValid;
  assign T83 = T77 ^ 1'h1;
  assign T84 = T80 ? 1'h1 : T85;
  assign T85 = T77 ? 1'h1 : 1'h0;
  assign T180 = T86[5'h1f:1'h0];
  assign T86 = T80 ? T89 : T87;
  assign T87 = T77 ? T88 : 38'h0;
  assign T88 = fifo_3_io_deqData[6'h25:1'h0];
  assign T89 = fifo_11_io_deqData[6'h25:1'h0];
  assign T90 = fifo_10_io_deqData[6'h2b:6'h26];
  assign T91 = fifo_2_io_deqData[6'h2b:6'h26];
  assign T92 = T98 ? T97 : T93;
  assign T93 = T95 ? T94 : 6'h0;
  assign T94 = fifo_2_io_deqData[6'h2b:6'h26];
  assign T95 = T96 & memoryBank_2_io_isWriteLoadRdy;
  assign T96 = fifo_2_io_deqValid;
  assign T97 = fifo_10_io_deqData[6'h2b:6'h26];
  assign T98 = T101 & T99;
  assign T99 = T100 & memoryBank_2_io_isWriteFabricRdy;
  assign T100 = fifo_10_io_deqValid;
  assign T101 = T95 ^ 1'h1;
  assign T102 = T98 ? 1'h1 : T103;
  assign T103 = T95 ? 1'h1 : 1'h0;
  assign T181 = T104[5'h1f:1'h0];
  assign T104 = T98 ? T107 : T105;
  assign T105 = T95 ? T106 : 38'h0;
  assign T106 = fifo_2_io_deqData[6'h25:1'h0];
  assign T107 = fifo_10_io_deqData[6'h25:1'h0];
  assign T108 = fifo_9_io_deqData[6'h2b:6'h26];
  assign T109 = fifo_1_io_deqData[6'h2b:6'h26];
  assign T110 = T116 ? T115 : T111;
  assign T111 = T113 ? T112 : 6'h0;
  assign T112 = fifo_1_io_deqData[6'h2b:6'h26];
  assign T113 = T114 & memoryBank_1_io_isWriteLoadRdy;
  assign T114 = fifo_1_io_deqValid;
  assign T115 = fifo_9_io_deqData[6'h2b:6'h26];
  assign T116 = T119 & T117;
  assign T117 = T118 & memoryBank_1_io_isWriteFabricRdy;
  assign T118 = fifo_9_io_deqValid;
  assign T119 = T113 ^ 1'h1;
  assign T120 = T116 ? 1'h1 : T121;
  assign T121 = T113 ? 1'h1 : 1'h0;
  assign T182 = T122[5'h1f:1'h0];
  assign T122 = T116 ? T125 : T123;
  assign T123 = T113 ? T124 : 38'h0;
  assign T124 = fifo_1_io_deqData[6'h25:1'h0];
  assign T125 = fifo_9_io_deqData[6'h25:1'h0];
  assign T126 = fifo_8_io_deqData[6'h2b:6'h26];
  assign T127 = fifo_io_deqData[6'h2b:6'h26];
  assign T128 = T134 ? T133 : T129;
  assign T129 = T131 ? T130 : 6'h0;
  assign T130 = fifo_io_deqData[6'h2b:6'h26];
  assign T131 = T132 & memoryBank_io_isWriteLoadRdy;
  assign T132 = fifo_io_deqValid;
  assign T133 = fifo_8_io_deqData[6'h2b:6'h26];
  assign T134 = T137 & T135;
  assign T135 = T136 & memoryBank_io_isWriteFabricRdy;
  assign T136 = fifo_8_io_deqValid;
  assign T137 = T131 ^ 1'h1;
  assign T138 = T134 ? 1'h1 : T139;
  assign T139 = T131 ? 1'h1 : 1'h0;
  assign T183 = T140[5'h1f:1'h0];
  assign T140 = T134 ? T143 : T141;
  assign T141 = T131 ? T142 : 38'h0;
  assign T142 = fifo_io_deqData[6'h25:1'h0];
  assign T143 = fifo_8_io_deqData[6'h25:1'h0];
  assign T144 = T8 ? memoryBank_7_io_isWriteFabricRdy : 1'h0;
  assign T184 = {6'h0, io_inDataFabric_7};
  assign T145 = T26 ? memoryBank_6_io_isWriteFabricRdy : 1'h0;
  assign T185 = {6'h0, io_inDataFabric_6};
  assign T146 = T44 ? memoryBank_5_io_isWriteFabricRdy : 1'h0;
  assign T186 = {6'h0, io_inDataFabric_5};
  assign T147 = T62 ? memoryBank_4_io_isWriteFabricRdy : 1'h0;
  assign T187 = {6'h0, io_inDataFabric_4};
  assign T148 = T80 ? memoryBank_3_io_isWriteFabricRdy : 1'h0;
  assign T188 = {6'h0, io_inDataFabric_3};
  assign T149 = T98 ? memoryBank_2_io_isWriteFabricRdy : 1'h0;
  assign T189 = {6'h0, io_inDataFabric_2};
  assign T150 = T116 ? memoryBank_1_io_isWriteFabricRdy : 1'h0;
  assign T190 = {6'h0, io_inDataFabric_1};
  assign T151 = T134 ? memoryBank_io_isWriteFabricRdy : 1'h0;
  assign T191 = {6'h0, io_inDataFabric_0};
  assign T152 = T5 ? memoryBank_7_io_isWriteLoadRdy : 1'h0;
  assign T192 = {6'h0, io_inDataLoad_7};
  assign T153 = T23 ? memoryBank_6_io_isWriteLoadRdy : 1'h0;
  assign T193 = {6'h0, io_inDataLoad_6};
  assign T154 = T41 ? memoryBank_5_io_isWriteLoadRdy : 1'h0;
  assign T194 = {6'h0, io_inDataLoad_5};
  assign T155 = T59 ? memoryBank_4_io_isWriteLoadRdy : 1'h0;
  assign T195 = {6'h0, io_inDataLoad_4};
  assign T156 = T77 ? memoryBank_3_io_isWriteLoadRdy : 1'h0;
  assign T196 = {6'h0, io_inDataLoad_3};
  assign T157 = T95 ? memoryBank_2_io_isWriteLoadRdy : 1'h0;
  assign T197 = {6'h0, io_inDataLoad_2};
  assign T158 = T113 ? memoryBank_1_io_isWriteLoadRdy : 1'h0;
  assign T198 = {6'h0, io_inDataLoad_1};
  assign T159 = T131 ? memoryBank_io_isWriteLoadRdy : 1'h0;
  assign T199 = {6'h0, io_inDataLoad_0};
  assign io_enqRdyFabric_0 = fifo_8_io_enqRdy;
  assign io_enqRdyFabric_1 = fifo_9_io_enqRdy;
  assign io_enqRdyFabric_2 = fifo_10_io_enqRdy;
  assign io_enqRdyFabric_3 = fifo_11_io_enqRdy;
  assign io_enqRdyFabric_4 = fifo_12_io_enqRdy;
  assign io_enqRdyFabric_5 = fifo_13_io_enqRdy;
  assign io_enqRdyFabric_6 = fifo_14_io_enqRdy;
  assign io_enqRdyFabric_7 = fifo_15_io_enqRdy;
  assign io_enqRdyLoad_0 = fifo_io_enqRdy;
  assign io_enqRdyLoad_1 = fifo_1_io_enqRdy;
  assign io_enqRdyLoad_2 = fifo_2_io_enqRdy;
  assign io_enqRdyLoad_3 = fifo_3_io_enqRdy;
  assign io_enqRdyLoad_4 = fifo_4_io_enqRdy;
  assign io_enqRdyLoad_5 = fifo_5_io_enqRdy;
  assign io_enqRdyLoad_6 = fifo_6_io_enqRdy;
  assign io_enqRdyLoad_7 = fifo_7_io_enqRdy;
  assign io_writeSuccess_0 = T160;
  assign T160 = T134 ? memoryBank_io_writeSuccess : T161;
  assign T161 = T131 ? memoryBank_io_writeSuccess : 1'h0;
  assign io_writeSuccess_1 = T162;
  assign T162 = T116 ? memoryBank_1_io_writeSuccess : T163;
  assign T163 = T113 ? memoryBank_1_io_writeSuccess : 1'h0;
  assign io_writeSuccess_2 = T164;
  assign T164 = T98 ? memoryBank_2_io_writeSuccess : T165;
  assign T165 = T95 ? memoryBank_2_io_writeSuccess : 1'h0;
  assign io_writeSuccess_3 = T166;
  assign T166 = T80 ? memoryBank_3_io_writeSuccess : T167;
  assign T167 = T77 ? memoryBank_3_io_writeSuccess : 1'h0;
  assign io_writeSuccess_4 = T168;
  assign T168 = T62 ? memoryBank_4_io_writeSuccess : T169;
  assign T169 = T59 ? memoryBank_4_io_writeSuccess : 1'h0;
  assign io_writeSuccess_5 = T170;
  assign T170 = T44 ? memoryBank_5_io_writeSuccess : T171;
  assign T171 = T41 ? memoryBank_5_io_writeSuccess : 1'h0;
  assign io_writeSuccess_6 = T172;
  assign T172 = T26 ? memoryBank_6_io_writeSuccess : T173;
  assign T173 = T23 ? memoryBank_6_io_writeSuccess : 1'h0;
  assign io_writeSuccess_7 = T174;
  assign T174 = T8 ? memoryBank_7_io_writeSuccess : T175;
  assign T175 = T5 ? memoryBank_7_io_writeSuccess : 1'h0;
  assign io_readSuccess_0 = memoryBank_io_readSuccess;
  assign io_readSuccess_1 = memoryBank_1_io_readSuccess;
  assign io_readSuccess_2 = memoryBank_2_io_readSuccess;
  assign io_readSuccess_3 = memoryBank_3_io_readSuccess;
  assign io_readSuccess_4 = memoryBank_4_io_readSuccess;
  assign io_readSuccess_5 = memoryBank_5_io_readSuccess;
  assign io_readSuccess_6 = memoryBank_6_io_readSuccess;
  assign io_readSuccess_7 = memoryBank_7_io_readSuccess;
  assign io_isReadValid_0 = memoryBank_io_isValid;
  assign io_isReadValid_1 = memoryBank_1_io_isValid;
  assign io_isReadValid_2 = memoryBank_2_io_isValid;
  assign io_isReadValid_3 = memoryBank_3_io_isValid;
  assign io_isReadValid_4 = memoryBank_4_io_isValid;
  assign io_isReadValid_5 = memoryBank_5_io_isValid;
  assign io_isReadValid_6 = memoryBank_6_io_isValid;
  assign io_isReadValid_7 = memoryBank_7_io_isValid;
  assign io_outData_0 = T200;
  assign T200 = {6'h0, memoryBank_io_outData};
  assign io_outData_1 = T201;
  assign T201 = {6'h0, memoryBank_1_io_outData};
  assign io_outData_2 = T202;
  assign T202 = {6'h0, memoryBank_2_io_outData};
  assign io_outData_3 = T203;
  assign T203 = {6'h0, memoryBank_3_io_outData};
  assign io_outData_4 = T204;
  assign T204 = {6'h0, memoryBank_4_io_outData};
  assign io_outData_5 = T205;
  assign T205 = {6'h0, memoryBank_5_io_outData};
  assign io_outData_6 = T206;
  assign T206 = {6'h0, memoryBank_6_io_outData};
  assign io_outData_7 = T207;
  assign T207 = {6'h0, memoryBank_7_io_outData};
  fifo_6 fifo(.clk(clk), .reset(reset),
       .io_enqData( T199 ),
       .io_deqData( fifo_io_deqData ),
       .io_enqRdy( fifo_io_enqRdy ),
       .io_deqRdy( T159 ),
       .io_enqValid( io_enqValidLoad_0 ),
       .io_deqValid( fifo_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_1(.clk(clk), .reset(reset),
       .io_enqData( T198 ),
       .io_deqData( fifo_1_io_deqData ),
       .io_enqRdy( fifo_1_io_enqRdy ),
       .io_deqRdy( T158 ),
       .io_enqValid( io_enqValidLoad_1 ),
       .io_deqValid( fifo_1_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_2(.clk(clk), .reset(reset),
       .io_enqData( T197 ),
       .io_deqData( fifo_2_io_deqData ),
       .io_enqRdy( fifo_2_io_enqRdy ),
       .io_deqRdy( T157 ),
       .io_enqValid( io_enqValidLoad_2 ),
       .io_deqValid( fifo_2_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_3(.clk(clk), .reset(reset),
       .io_enqData( T196 ),
       .io_deqData( fifo_3_io_deqData ),
       .io_enqRdy( fifo_3_io_enqRdy ),
       .io_deqRdy( T156 ),
       .io_enqValid( io_enqValidLoad_3 ),
       .io_deqValid( fifo_3_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_4(.clk(clk), .reset(reset),
       .io_enqData( T195 ),
       .io_deqData( fifo_4_io_deqData ),
       .io_enqRdy( fifo_4_io_enqRdy ),
       .io_deqRdy( T155 ),
       .io_enqValid( io_enqValidLoad_4 ),
       .io_deqValid( fifo_4_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_5(.clk(clk), .reset(reset),
       .io_enqData( T194 ),
       .io_deqData( fifo_5_io_deqData ),
       .io_enqRdy( fifo_5_io_enqRdy ),
       .io_deqRdy( T154 ),
       .io_enqValid( io_enqValidLoad_5 ),
       .io_deqValid( fifo_5_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_6(.clk(clk), .reset(reset),
       .io_enqData( T193 ),
       .io_deqData( fifo_6_io_deqData ),
       .io_enqRdy( fifo_6_io_enqRdy ),
       .io_deqRdy( T153 ),
       .io_enqValid( io_enqValidLoad_6 ),
       .io_deqValid( fifo_6_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_7(.clk(clk), .reset(reset),
       .io_enqData( T192 ),
       .io_deqData( fifo_7_io_deqData ),
       .io_enqRdy( fifo_7_io_enqRdy ),
       .io_deqRdy( T152 ),
       .io_enqValid( io_enqValidLoad_7 ),
       .io_deqValid( fifo_7_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_8(.clk(clk), .reset(reset),
       .io_enqData( T191 ),
       .io_deqData( fifo_8_io_deqData ),
       .io_enqRdy( fifo_8_io_enqRdy ),
       .io_deqRdy( T151 ),
       .io_enqValid( io_enqValidFabric_0 ),
       .io_deqValid( fifo_8_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_9(.clk(clk), .reset(reset),
       .io_enqData( T190 ),
       .io_deqData( fifo_9_io_deqData ),
       .io_enqRdy( fifo_9_io_enqRdy ),
       .io_deqRdy( T150 ),
       .io_enqValid( io_enqValidFabric_1 ),
       .io_deqValid( fifo_9_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_10(.clk(clk), .reset(reset),
       .io_enqData( T189 ),
       .io_deqData( fifo_10_io_deqData ),
       .io_enqRdy( fifo_10_io_enqRdy ),
       .io_deqRdy( T149 ),
       .io_enqValid( io_enqValidFabric_2 ),
       .io_deqValid( fifo_10_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_11(.clk(clk), .reset(reset),
       .io_enqData( T188 ),
       .io_deqData( fifo_11_io_deqData ),
       .io_enqRdy( fifo_11_io_enqRdy ),
       .io_deqRdy( T148 ),
       .io_enqValid( io_enqValidFabric_3 ),
       .io_deqValid( fifo_11_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_12(.clk(clk), .reset(reset),
       .io_enqData( T187 ),
       .io_deqData( fifo_12_io_deqData ),
       .io_enqRdy( fifo_12_io_enqRdy ),
       .io_deqRdy( T147 ),
       .io_enqValid( io_enqValidFabric_4 ),
       .io_deqValid( fifo_12_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_13(.clk(clk), .reset(reset),
       .io_enqData( T186 ),
       .io_deqData( fifo_13_io_deqData ),
       .io_enqRdy( fifo_13_io_enqRdy ),
       .io_deqRdy( T146 ),
       .io_enqValid( io_enqValidFabric_5 ),
       .io_deqValid( fifo_13_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_14(.clk(clk), .reset(reset),
       .io_enqData( T185 ),
       .io_deqData( fifo_14_io_deqData ),
       .io_enqRdy( fifo_14_io_enqRdy ),
       .io_deqRdy( T145 ),
       .io_enqValid( io_enqValidFabric_6 ),
       .io_deqValid( fifo_14_io_deqValid ),
       .io_rst( io_rst )
  );
  fifo_6 fifo_15(.clk(clk), .reset(reset),
       .io_enqData( T184 ),
       .io_deqData( fifo_15_io_deqData ),
       .io_enqRdy( fifo_15_io_enqRdy ),
       .io_deqRdy( T144 ),
       .io_enqValid( io_enqValidFabric_7 ),
       .io_deqValid( fifo_15_io_deqValid ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank(.clk(clk), .reset(reset),
       .io_inData( T183 ),
       .io_outData( memoryBank_io_outData ),
       .io_readEn( io_readEn_0 ),
       .io_writeEn( T138 ),
       .io_writeSuccess( memoryBank_io_writeSuccess ),
       .io_readSuccess( memoryBank_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_0 ),
       .io_isValid( memoryBank_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_0 ),
       .io_writeAddr( T128 ),
       .io_writeLoadAddr( T127 ),
       .io_writeFabricAddr( T126 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_1(.clk(clk), .reset(reset),
       .io_inData( T182 ),
       .io_outData( memoryBank_1_io_outData ),
       .io_readEn( io_readEn_1 ),
       .io_writeEn( T120 ),
       .io_writeSuccess( memoryBank_1_io_writeSuccess ),
       .io_readSuccess( memoryBank_1_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_1 ),
       .io_isValid( memoryBank_1_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_1_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_1_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_1 ),
       .io_writeAddr( T110 ),
       .io_writeLoadAddr( T109 ),
       .io_writeFabricAddr( T108 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_2(.clk(clk), .reset(reset),
       .io_inData( T181 ),
       .io_outData( memoryBank_2_io_outData ),
       .io_readEn( io_readEn_2 ),
       .io_writeEn( T102 ),
       .io_writeSuccess( memoryBank_2_io_writeSuccess ),
       .io_readSuccess( memoryBank_2_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_2 ),
       .io_isValid( memoryBank_2_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_2_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_2_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_2 ),
       .io_writeAddr( T92 ),
       .io_writeLoadAddr( T91 ),
       .io_writeFabricAddr( T90 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_3(.clk(clk), .reset(reset),
       .io_inData( T180 ),
       .io_outData( memoryBank_3_io_outData ),
       .io_readEn( io_readEn_3 ),
       .io_writeEn( T84 ),
       .io_writeSuccess( memoryBank_3_io_writeSuccess ),
       .io_readSuccess( memoryBank_3_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_3 ),
       .io_isValid( memoryBank_3_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_3_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_3_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_3 ),
       .io_writeAddr( T74 ),
       .io_writeLoadAddr( T73 ),
       .io_writeFabricAddr( T72 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_4(.clk(clk), .reset(reset),
       .io_inData( T179 ),
       .io_outData( memoryBank_4_io_outData ),
       .io_readEn( io_readEn_4 ),
       .io_writeEn( T66 ),
       .io_writeSuccess( memoryBank_4_io_writeSuccess ),
       .io_readSuccess( memoryBank_4_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_4 ),
       .io_isValid( memoryBank_4_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_4_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_4_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_4 ),
       .io_writeAddr( T56 ),
       .io_writeLoadAddr( T55 ),
       .io_writeFabricAddr( T54 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_5(.clk(clk), .reset(reset),
       .io_inData( T178 ),
       .io_outData( memoryBank_5_io_outData ),
       .io_readEn( io_readEn_5 ),
       .io_writeEn( T48 ),
       .io_writeSuccess( memoryBank_5_io_writeSuccess ),
       .io_readSuccess( memoryBank_5_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_5 ),
       .io_isValid( memoryBank_5_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_5_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_5_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_5 ),
       .io_writeAddr( T38 ),
       .io_writeLoadAddr( T37 ),
       .io_writeFabricAddr( T36 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_6(.clk(clk), .reset(reset),
       .io_inData( T177 ),
       .io_outData( memoryBank_6_io_outData ),
       .io_readEn( io_readEn_6 ),
       .io_writeEn( T30 ),
       .io_writeSuccess( memoryBank_6_io_writeSuccess ),
       .io_readSuccess( memoryBank_6_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_6 ),
       .io_isValid( memoryBank_6_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_6_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_6_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_6 ),
       .io_writeAddr( T20 ),
       .io_writeLoadAddr( T19 ),
       .io_writeFabricAddr( T18 ),
       .io_rst( io_rst )
  );
  memoryBank memoryBank_7(.clk(clk), .reset(reset),
       .io_inData( T176 ),
       .io_outData( memoryBank_7_io_outData ),
       .io_readEn( io_readEn_7 ),
       .io_writeEn( T12 ),
       .io_writeSuccess( memoryBank_7_io_writeSuccess ),
       .io_readSuccess( memoryBank_7_io_readSuccess ),
       .io_doInvalidate( io_doInvalidate_7 ),
       .io_isValid( memoryBank_7_io_isValid ),
       .io_isWriteLoadRdy( memoryBank_7_io_isWriteLoadRdy ),
       .io_isWriteFabricRdy( memoryBank_7_io_isWriteFabricRdy ),
       .io_readAddr( io_readAddr_7 ),
       .io_writeAddr( T2 ),
       .io_writeLoadAddr( T1 ),
       .io_writeFabricAddr( T0 ),
       .io_rst( io_rst )
  );
endmodule

module memConfig_0(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[8:0] io_memAddr,
    output[88:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T94;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T95;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T96;
  reg  iterCnt;
  wire T97;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T98;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T99;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[88:0] T100;
  wire[92:0] T76;
  wire[92:0] T77;
  wire[61:0] T78;
  reg [30:0] memData_0;
  wire[30:0] T101;
  wire[30:0] T79;
  wire[30:0] T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  wire[1:0] T84;
  wire[1:0] T102;
  reg [30:0] memData_1;
  wire[30:0] T103;
  wire[30:0] T85;
  wire T86;
  wire T87;
  reg [30:0] memData_2;
  wire[30:0] T104;
  wire[30:0] T88;
  wire T89;
  wire T90;
  wire[8:0] T91;
  reg [8:0] memAddr;
  wire[8:0] T105;
  wire[8:0] T92;
  wire[8:0] T93;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memData_2 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T94 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T95 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = T96 == 2'h2;
  assign T96 = {1'h0, iterCnt};
  assign T97 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = T98 < 2'h2;
  assign T98 = {1'h0, iterCnt};
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T99 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'hc;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'hc;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'hc;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'hc;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T100;
  assign T100 = T76[7'h58:1'h0];
  assign T76 = memOutValid ? T77 : 93'h0;
  assign T77 = {memData_2, T78};
  assign T78 = {memData_1, memData_0};
  assign T101 = reset ? 31'h0 : T79;
  assign T79 = T81 ? T80 : memData_0;
  assign T80 = inConfigReg[5'h1e:1'h0];
  assign T81 = T45 & T82;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = 1'h1 << T84;
  assign T84 = T102;
  assign T102 = {1'h0, iterCnt};
  assign T103 = reset ? 31'h0 : T85;
  assign T85 = T86 ? T80 : memData_1;
  assign T86 = T45 & T87;
  assign T87 = T83[1'h1:1'h1];
  assign T104 = reset ? 31'h0 : T88;
  assign T88 = T89 ? T80 : memData_2;
  assign T89 = T45 & T90;
  assign T90 = T83[2'h2:2'h2];
  assign io_memAddr = T91;
  assign T91 = memOutValid ? memAddr : 9'h0;
  assign T105 = reset ? 9'h0 : T92;
  assign T92 = memOutValid ? T93 : memAddr;
  assign T93 = memAddr + 9'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T81) begin
      memData_0 <= T80;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T86) begin
      memData_1 <= T80;
    end
    if(reset) begin
      memData_2 <= 31'h0;
    end else if(T89) begin
      memData_2 <= T80;
    end
    if(reset) begin
      memAddr <= 9'h0;
    end else if(memOutValid) begin
      memAddr <= T93;
    end
  end
endmodule

module fifo_0(input clk, input reset,
    input [31:0] io_enqData,
    output[31:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg [1:0] deqPtr;
  wire[1:0] T21;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] deqPtrInc;
  wire[1:0] T4;
  wire doDeq;
  wire T5;
  reg [1:0] enqPtr;
  wire[1:0] T22;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] enqPtrInc;
  wire[1:0] T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[31:0] T19;
  reg [31:0] fifoMem [3:0];
  wire[31:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      fifoMem[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 2'h0 : T2;
  assign T2 = io_rst ? 2'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 3'h4;
  assign T4 = deqPtr + 2'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 2'h0 : T6;
  assign T6 = io_rst ? 2'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 3'h4;
  assign T8 = enqPtr + 2'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 2'h0;
    end else if(io_rst) begin
      deqPtr <= 2'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 2'h0;
    end else if(io_rst) begin
      enqPtr <= 2'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fifo_1(input clk, input reset,
    input [31:0] io_enqData,
    output[31:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg  deqPtr;
  wire T21;
  wire T2;
  wire T3;
  wire deqPtrInc;
  wire T4;
  wire doDeq;
  wire T5;
  reg  enqPtr;
  wire T22;
  wire T6;
  wire T7;
  wire enqPtrInc;
  wire T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[31:0] T19;
  reg [31:0] fifoMem [1:0];
  wire[31:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      fifoMem[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = io_rst ? 1'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 2'h2;
  assign T4 = deqPtr + 1'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 1'h0 : T6;
  assign T6 = io_rst ? 1'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 2'h2;
  assign T8 = enqPtr + 1'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(io_rst) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(io_rst) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fabInSeqDP(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input [8:0] io_seqMemAddr,
    input  io_seqMemAddrValid,
    output[31:0] io_fabInData_19,
    output[31:0] io_fabInData_18,
    output[31:0] io_fabInData_17,
    output[31:0] io_fabInData_16,
    output[31:0] io_fabInData_15,
    output[31:0] io_fabInData_14,
    output[31:0] io_fabInData_13,
    output[31:0] io_fabInData_12,
    output[31:0] io_fabInData_11,
    output[31:0] io_fabInData_10,
    output[31:0] io_fabInData_9,
    output[31:0] io_fabInData_8,
    output[31:0] io_fabInData_7,
    output[31:0] io_fabInData_6,
    output[31:0] io_fabInData_5,
    output[31:0] io_fabInData_4,
    output[31:0] io_fabInData_3,
    output[31:0] io_fabInData_2,
    output[31:0] io_fabInData_1,
    output[31:0] io_fabInData_0,
    output io_fabInValid_19,
    output io_fabInValid_18,
    output io_fabInValid_17,
    output io_fabInValid_16,
    output io_fabInValid_15,
    output io_fabInValid_14,
    output io_fabInValid_13,
    output io_fabInValid_12,
    output io_fabInValid_11,
    output io_fabInValid_10,
    output io_fabInValid_9,
    output io_fabInValid_8,
    output io_fabInValid_7,
    output io_fabInValid_6,
    output io_fabInValid_5,
    output io_fabInValid_4,
    output io_fabInValid_3,
    output io_fabInValid_2,
    output io_fabInValid_1,
    output io_fabInValid_0,
    input  io_fabInRdy_19,
    input  io_fabInRdy_18,
    input  io_fabInRdy_17,
    input  io_fabInRdy_16,
    input  io_fabInRdy_15,
    input  io_fabInRdy_14,
    input  io_fabInRdy_13,
    input  io_fabInRdy_12,
    input  io_fabInRdy_11,
    input  io_fabInRdy_10,
    input  io_fabInRdy_9,
    input  io_fabInRdy_8,
    input  io_fabInRdy_7,
    input  io_fabInRdy_6,
    input  io_fabInRdy_5,
    input  io_fabInRdy_4,
    input  io_fabInRdy_3,
    input  io_fabInRdy_2,
    input  io_fabInRdy_1,
    input  io_fabInRdy_0,
    input [37:0] io_loadStore_7,
    input [37:0] io_loadStore_6,
    input [37:0] io_loadStore_5,
    input [37:0] io_loadStore_4,
    input [37:0] io_loadStore_3,
    input [37:0] io_loadStore_2,
    input [37:0] io_loadStore_1,
    input [37:0] io_loadStore_0,
    input  io_loadStoreValid_7,
    input  io_loadStoreValid_6,
    input  io_loadStoreValid_5,
    input  io_loadStoreValid_4,
    input  io_loadStoreValid_3,
    input  io_loadStoreValid_2,
    input  io_loadStoreValid_1,
    input  io_loadStoreValid_0,
    output io_loadStoreRdy_7,
    output io_loadStoreRdy_6,
    output io_loadStoreRdy_5,
    output io_loadStoreRdy_4,
    output io_loadStoreRdy_3,
    output io_loadStoreRdy_2,
    output io_loadStoreRdy_1,
    output io_loadStoreRdy_0,
    input [37:0] io_fabStore_7,
    input [37:0] io_fabStore_6,
    input [37:0] io_fabStore_5,
    input [37:0] io_fabStore_4,
    input [37:0] io_fabStore_3,
    input [37:0] io_fabStore_2,
    input [37:0] io_fabStore_1,
    input [37:0] io_fabStore_0,
    input  io_fabStoreValid_7,
    input  io_fabStoreValid_6,
    input  io_fabStoreValid_5,
    input  io_fabStoreValid_4,
    input  io_fabStoreValid_3,
    input  io_fabStoreValid_2,
    input  io_fabStoreValid_1,
    input  io_fabStoreValid_0,
    output io_fabStoreRdy_7,
    output io_fabStoreRdy_6,
    output io_fabStoreRdy_5,
    output io_fabStoreRdy_4,
    output io_fabStoreRdy_3,
    output io_fabStoreRdy_2,
    output io_fabStoreRdy_1,
    output io_fabStoreRdy_0,
    output io_seqProceed
);

  wire T0;
  wire T1;
  wire isReadValid;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[87:0] bankSeq;
  wire[87:0] T20;
  wire[87:0] T21;
  wire[87:0] T22;
  wire[87:0] T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[87:0] T26;
  wire[87:0] T27;
  wire[87:0] T28;
  wire[87:0] T29;
  wire[87:0] T30;
  wire[87:0] T31;
  wire[87:0] T32;
  wire[87:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[88:0] nextSeq;
  wire[88:0] T36;
  wire[88:0] T37;
  wire[88:0] T38;
  wire[88:0] T39;
  wire[88:0] T40;
  wire[88:0] T41;
  wire[88:0] T42;
  wire[88:0] T43;
  wire[88:0] T44;
  wire[88:0] T45;
  wire[88:0] T46;
  wire[88:0] T47;
  wire[88:0] T48;
  wire[88:0] T49;
  wire[88:0] T50;
  wire[88:0] T51;
  wire[88:0] T52;
  wire[88:0] T53;
  wire[88:0] T54;
  wire[88:0] T55;
  wire[88:0] T56;
  wire[88:0] T57;
  wire[88:0] T58;
  wire T59;
  reg  nextSeqSelReg;
  wire T3098;
  wire T60;
  wire T61;
  wire T62;
  wire allDone;
  wire T63;
  wire bankReadDone_7;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire bankReadDone_6;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire bankReadDone_5;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire bankReadDone_4;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire bankReadDone_3;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire bankReadDone_2;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire bankReadDone_1;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire bankReadDone_0;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  reg [88:0] nextSeqReg2;
  wire[88:0] T3099;
  wire[88:0] T170;
  wire[88:0] nextSeqWire;
  wire[88:0] T171;
  wire[88:0] T172;
  wire T173;
  wire T174;
  reg  firstSeqSelReg;
  wire T3100;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[87:0] T182;
  wire T183;
  reg  bankReadDoneReg_1;
  wire T3101;
  wire T184;
  wire readDone_1;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  reg  nextSeqRegValid2;
  wire T3102;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  reg  nextSeqRegValid1;
  wire T3103;
  wire T197;
  wire T198;
  wire[87:0] T199;
  wire T200;
  reg  bankReadDoneReg_2;
  wire T3104;
  wire T201;
  wire readDone_2;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire[87:0] T207;
  wire T208;
  reg  bankReadDoneReg_3;
  wire T3105;
  wire T209;
  wire readDone_3;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[87:0] T215;
  wire T216;
  reg  bankReadDoneReg_4;
  wire T3106;
  wire T217;
  wire readDone_4;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire[87:0] T223;
  wire T224;
  reg  bankReadDoneReg_5;
  wire T3107;
  wire T225;
  wire readDone_5;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[87:0] T231;
  wire T232;
  reg  bankReadDoneReg_6;
  wire T3108;
  wire T233;
  wire readDone_6;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire[87:0] T239;
  wire T240;
  reg  bankReadDoneReg_7;
  wire T3109;
  wire T241;
  wire readDone_7;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  reg  bankReadDoneReg_0;
  wire T3110;
  wire T248;
  wire readDone_0;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire collectRdy;
  wire T270;
  wire T271;
  wire T272;
  wire rdy;
  wire T273;
  wire T274;
  wire T275;
  wire enqRdyCollect_19;
  wire T276;
  wire T277;
  wire enqRdyCollect_18;
  wire T278;
  wire T279;
  wire enqRdyCollect_17;
  wire T280;
  wire T281;
  wire enqRdyCollect_16;
  wire T282;
  wire T283;
  wire enqRdyCollect_15;
  wire T284;
  wire T285;
  wire enqRdyCollect_14;
  wire T286;
  wire T287;
  wire enqRdyCollect_13;
  wire T288;
  wire T289;
  wire enqRdyCollect_12;
  wire T290;
  wire T291;
  wire enqRdyCollect_11;
  wire T292;
  wire T293;
  wire enqRdyCollect_10;
  wire T294;
  wire T295;
  wire enqRdyCollect_9;
  wire T296;
  wire T297;
  wire enqRdyCollect_8;
  wire T298;
  wire T299;
  wire enqRdyCollect_7;
  wire T300;
  wire T301;
  wire enqRdyCollect_6;
  wire T302;
  wire T303;
  wire enqRdyCollect_5;
  wire T304;
  wire T305;
  wire enqRdyCollect_4;
  wire T306;
  wire T307;
  wire enqRdyCollect_3;
  wire T308;
  wire T309;
  wire enqRdyCollect_2;
  wire T310;
  wire T311;
  wire enqRdyCollect_1;
  wire T312;
  wire enqRdyCollect_0;
  wire T313;
  wire rdyInit;
  wire T314;
  reg  seqLevelDoneReg2;
  wire T3111;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T361;
  wire T362;
  wire T363;
  wire bankToPortValid_7_0;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[31:0] T368;
  wire[4:0] T369;
  wire[4:0] T3112;
  wire[2:0] portId;
  wire[2:0] T370;
  wire[2:0] T371;
  wire[2:0] T372;
  wire[2:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire[2:0] T376;
  wire[2:0] T377;
  wire[2:0] T378;
  wire[2:0] T379;
  wire[2:0] T380;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire[87:0] bankSeq2;
  wire[87:0] T386;
  wire[87:0] T387;
  wire[87:0] T388;
  wire[87:0] T389;
  wire[87:0] T390;
  wire[87:0] T391;
  wire[87:0] T392;
  wire[87:0] T393;
  wire[87:0] T394;
  wire[87:0] T395;
  wire[87:0] T396;
  wire[87:0] T397;
  wire[87:0] T398;
  wire[87:0] T399;
  wire[87:0] T400;
  reg [87:0] bankSeqReg_0;
  wire[87:0] T3113;
  reg [87:0] bankSeqReg_1;
  wire[87:0] T3114;
  reg [87:0] bankSeqReg_2;
  wire[87:0] T3115;
  reg [87:0] bankSeqReg_3;
  wire[87:0] T3116;
  reg [87:0] bankSeqReg_4;
  wire[87:0] T3117;
  reg [87:0] bankSeqReg_5;
  wire[87:0] T3118;
  reg [87:0] bankSeqReg_6;
  wire[87:0] T3119;
  reg [87:0] bankSeqReg_7;
  wire[87:0] T3120;
  wire[2:0] T401;
  wire T402;
  wire T403;
  wire[2:0] T404;
  wire T405;
  wire T406;
  wire[2:0] T407;
  wire T408;
  wire[2:0] T409;
  wire T410;
  wire T411;
  wire[2:0] T412;
  wire T413;
  wire[2:0] T414;
  wire T415;
  wire T416;
  wire[2:0] T417;
  wire T418;
  wire[2:0] T419;
  wire T420;
  wire T421;
  wire[2:0] T422;
  wire T423;
  wire[2:0] T424;
  wire T425;
  wire T426;
  wire[2:0] T427;
  wire T428;
  wire[2:0] T429;
  wire T430;
  wire T431;
  wire[2:0] T432;
  wire T433;
  wire[2:0] T434;
  wire[2:0] T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire bankToPortValid_6_0;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[31:0] T444;
  wire[4:0] T445;
  wire[4:0] T3121;
  wire T446;
  wire T447;
  wire T448;
  wire bankToPortValid_5_0;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire[31:0] T453;
  wire[4:0] T454;
  wire[4:0] T3122;
  wire T455;
  wire T456;
  wire T457;
  wire bankToPortValid_4_0;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire[31:0] T462;
  wire[4:0] T463;
  wire[4:0] T3123;
  wire T464;
  wire T465;
  wire T466;
  wire bankToPortValid_3_0;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[31:0] T471;
  wire[4:0] T472;
  wire[4:0] T3124;
  wire T473;
  wire T474;
  wire T475;
  wire bankToPortValid_2_0;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire[31:0] T480;
  wire[4:0] T481;
  wire[4:0] T3125;
  wire T482;
  wire T483;
  wire T484;
  wire bankToPortValid_1_0;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire[31:0] T489;
  wire[4:0] T490;
  wire[4:0] T3126;
  wire T491;
  wire T492;
  wire bankToPortValid_0_0;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire[31:0] T497;
  wire[4:0] T498;
  wire[4:0] T3127;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire bankToPortValid_7_1;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire bankToPortValid_6_1;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire bankToPortValid_5_1;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire bankToPortValid_4_1;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire bankToPortValid_3_1;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire bankToPortValid_2_1;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire bankToPortValid_1_1;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire bankToPortValid_0_1;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire bankToPortValid_7_2;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire bankToPortValid_6_2;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire bankToPortValid_5_2;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire bankToPortValid_4_2;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire bankToPortValid_3_2;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire bankToPortValid_2_2;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire bankToPortValid_1_2;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire bankToPortValid_0_2;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire bankToPortValid_7_3;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire bankToPortValid_6_3;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire bankToPortValid_5_3;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire bankToPortValid_4_3;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire bankToPortValid_3_3;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire bankToPortValid_2_3;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire bankToPortValid_1_3;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire bankToPortValid_0_3;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire bankToPortValid_7_4;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire bankToPortValid_6_4;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire bankToPortValid_5_4;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire bankToPortValid_4_4;
  wire T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire bankToPortValid_3_4;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire bankToPortValid_2_4;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire bankToPortValid_1_4;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire bankToPortValid_0_4;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire bankToPortValid_7_5;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire bankToPortValid_6_5;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire bankToPortValid_5_5;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire bankToPortValid_4_5;
  wire T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire bankToPortValid_3_5;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire bankToPortValid_2_5;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire bankToPortValid_1_5;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire bankToPortValid_0_5;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire bankToPortValid_7_6;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire bankToPortValid_6_6;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire bankToPortValid_5_6;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire bankToPortValid_4_6;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire bankToPortValid_3_6;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire bankToPortValid_2_6;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire bankToPortValid_1_6;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire bankToPortValid_0_6;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire bankToPortValid_7_7;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire bankToPortValid_6_7;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire bankToPortValid_5_7;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire bankToPortValid_4_7;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire bankToPortValid_3_7;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire bankToPortValid_2_7;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire bankToPortValid_1_7;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire bankToPortValid_0_7;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire bankToPortValid_7_8;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire T902;
  wire bankToPortValid_6_8;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire bankToPortValid_5_8;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire bankToPortValid_4_8;
  wire T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire bankToPortValid_3_8;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire bankToPortValid_2_8;
  wire T931;
  wire T932;
  wire T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire bankToPortValid_1_8;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire bankToPortValid_0_8;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire bankToPortValid_7_9;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire bankToPortValid_6_9;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire bankToPortValid_5_9;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire bankToPortValid_4_9;
  wire T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire bankToPortValid_3_9;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire bankToPortValid_2_9;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire bankToPortValid_1_9;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire bankToPortValid_0_9;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire T1006;
  wire T1007;
  wire bankToPortValid_7_10;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire bankToPortValid_6_10;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire bankToPortValid_5_10;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire bankToPortValid_4_10;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire bankToPortValid_3_10;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire bankToPortValid_2_10;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire bankToPortValid_1_10;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire T1055;
  wire bankToPortValid_0_10;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire bankToPortValid_7_11;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire bankToPortValid_6_11;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire bankToPortValid_5_11;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire bankToPortValid_4_11;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire bankToPortValid_3_11;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire bankToPortValid_2_11;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire bankToPortValid_1_11;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire bankToPortValid_0_11;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire bankToPortValid_7_12;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire bankToPortValid_6_12;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire T1133;
  wire bankToPortValid_5_12;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire bankToPortValid_4_12;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire bankToPortValid_3_12;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire bankToPortValid_2_12;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire bankToPortValid_1_12;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire bankToPortValid_0_12;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire bankToPortValid_7_13;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire bankToPortValid_6_13;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire bankToPortValid_5_13;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire bankToPortValid_4_13;
  wire T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire bankToPortValid_3_13;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire bankToPortValid_2_13;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire bankToPortValid_1_13;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire bankToPortValid_0_13;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire bankToPortValid_7_14;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire bankToPortValid_6_14;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire bankToPortValid_5_14;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire bankToPortValid_4_14;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire bankToPortValid_3_14;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire bankToPortValid_2_14;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire bankToPortValid_1_14;
  wire T1274;
  wire T1275;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire bankToPortValid_0_14;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire bankToPortValid_7_15;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  wire T1294;
  wire bankToPortValid_6_15;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire bankToPortValid_5_15;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire bankToPortValid_4_15;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire bankToPortValid_3_15;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire bankToPortValid_2_15;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire bankToPortValid_1_15;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire bankToPortValid_0_15;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire T1343;
  wire bankToPortValid_7_16;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire bankToPortValid_6_16;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire bankToPortValid_5_16;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire bankToPortValid_4_16;
  wire T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire bankToPortValid_3_16;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire bankToPortValid_2_16;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire bankToPortValid_1_16;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire bankToPortValid_0_16;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire bankToPortValid_7_17;
  wire T1400;
  wire T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire bankToPortValid_6_17;
  wire T1407;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire bankToPortValid_5_17;
  wire T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire bankToPortValid_4_17;
  wire T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire bankToPortValid_3_17;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire bankToPortValid_2_17;
  wire T1435;
  wire T1436;
  wire T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire bankToPortValid_1_17;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire bankToPortValid_0_17;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire bankToPortValid_7_18;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire bankToPortValid_6_18;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire bankToPortValid_5_18;
  wire T1470;
  wire T1471;
  wire T1472;
  wire T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire bankToPortValid_4_18;
  wire T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire bankToPortValid_3_18;
  wire T1484;
  wire T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire bankToPortValid_2_18;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire T1497;
  wire bankToPortValid_1_18;
  wire T1498;
  wire T1499;
  wire T1500;
  wire T1501;
  wire T1502;
  wire T1503;
  wire bankToPortValid_0_18;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire T1508;
  reg  seqLevelDoneReg1;
  wire T3128;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T1509;
  wire T1510;
  wire T1511;
  wire bankToPortValid_7_19;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire T1516;
  wire T1517;
  wire T1518;
  wire bankToPortValid_6_19;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire bankToPortValid_5_19;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire T1532;
  wire bankToPortValid_4_19;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire bankToPortValid_3_19;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  wire T1546;
  wire bankToPortValid_2_19;
  wire T1547;
  wire T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire T1553;
  wire bankToPortValid_1_19;
  wire T1554;
  wire T1555;
  wire T1556;
  wire T1557;
  wire T1558;
  wire T1559;
  wire bankToPortValid_0_19;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[31:0] T1569;
  wire[31:0] readValuelocStrg;
  wire[31:0] T3129;
  wire[37:0] T1570;
  wire[37:0] T1571;
  wire[37:0] T1572;
  wire[37:0] T1573;
  wire[37:0] T1574;
  wire[37:0] T1575;
  wire[37:0] T1576;
  wire[37:0] T1577;
  wire[37:0] T1578;
  wire[37:0] T1579;
  wire[37:0] T1580;
  wire[37:0] T1581;
  wire[37:0] T1582;
  wire[37:0] T1583;
  wire[37:0] T1584;
  wire T1585;
  wire T1586;
  wire T1587;
  wire[31:0] T1588;
  wire T1589;
  wire T1590;
  wire T1591;
  wire[31:0] T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire[31:0] T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire[31:0] T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire[31:0] T1604;
  wire T1605;
  wire T1606;
  wire T1607;
  wire[31:0] T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[31:0] T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[31:0] T1617;
  wire[31:0] T1618;
  wire[31:0] T1619;
  wire[31:0] T1620;
  wire[31:0] T1621;
  wire[31:0] T1622;
  wire[31:0] bankToPort_7_19;
  wire[31:0] T1623;
  wire[31:0] T1624;
  wire T1625;
  wire T1626;
  wire[31:0] T1627;
  wire[4:0] T1628;
  wire[4:0] T3130;
  wire[31:0] readValueBankFifo;
  wire[31:0] T1629;
  wire[31:0] T1630;
  wire[31:0] T1631;
  wire[31:0] T1632;
  wire[31:0] T1633;
  wire[31:0] T1634;
  wire[31:0] T1635;
  wire[31:0] T1636;
  wire[31:0] T1637;
  wire[31:0] T1638;
  wire[31:0] T1639;
  wire[31:0] T1640;
  wire[31:0] T1641;
  wire[31:0] T1642;
  wire[31:0] T1643;
  wire T1644;
  wire[31:0] T1645;
  wire[31:0] T1646;
  wire[31:0] bankToPort_6_19;
  wire[31:0] T1647;
  wire[31:0] T1648;
  wire T1649;
  wire T1650;
  wire[31:0] T1651;
  wire[4:0] T1652;
  wire[4:0] T3131;
  wire T1653;
  wire[31:0] T1654;
  wire[31:0] T1655;
  wire[31:0] bankToPort_5_19;
  wire[31:0] T1656;
  wire[31:0] T1657;
  wire T1658;
  wire T1659;
  wire[31:0] T1660;
  wire[4:0] T1661;
  wire[4:0] T3132;
  wire T1662;
  wire[31:0] T1663;
  wire[31:0] T1664;
  wire[31:0] bankToPort_4_19;
  wire[31:0] T1665;
  wire[31:0] T1666;
  wire T1667;
  wire T1668;
  wire[31:0] T1669;
  wire[4:0] T1670;
  wire[4:0] T3133;
  wire T1671;
  wire[31:0] T1672;
  wire[31:0] T1673;
  wire[31:0] bankToPort_3_19;
  wire[31:0] T1674;
  wire[31:0] T1675;
  wire T1676;
  wire T1677;
  wire[31:0] T1678;
  wire[4:0] T1679;
  wire[4:0] T3134;
  wire T1680;
  wire[31:0] T1681;
  wire[31:0] T1682;
  wire[31:0] bankToPort_2_19;
  wire[31:0] T1683;
  wire[31:0] T1684;
  wire T1685;
  wire T1686;
  wire[31:0] T1687;
  wire[4:0] T1688;
  wire[4:0] T3135;
  wire T1689;
  wire[31:0] T1690;
  wire[31:0] T1691;
  wire[31:0] bankToPort_1_19;
  wire[31:0] T1692;
  wire[31:0] T1693;
  wire T1694;
  wire T1695;
  wire[31:0] T1696;
  wire[4:0] T1697;
  wire[4:0] T3136;
  wire T1698;
  wire[31:0] T1699;
  wire[31:0] T1700;
  wire[31:0] bankToPort_0_19;
  wire[31:0] T1701;
  wire[31:0] T1702;
  wire T1703;
  wire T1704;
  wire[31:0] T1705;
  wire[4:0] T1706;
  wire[4:0] T3137;
  wire T1707;
  wire T1708;
  wire T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[31:0] T1713;
  wire[31:0] T1714;
  wire[31:0] T1715;
  wire[31:0] T1716;
  wire[31:0] T1717;
  wire[31:0] T1718;
  wire[31:0] bankToPort_7_18;
  wire[31:0] T1719;
  wire[31:0] T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[31:0] T1724;
  wire[31:0] T1725;
  wire[31:0] bankToPort_6_18;
  wire[31:0] T1726;
  wire[31:0] T1727;
  wire T1728;
  wire T1729;
  wire T1730;
  wire[31:0] T1731;
  wire[31:0] T1732;
  wire[31:0] bankToPort_5_18;
  wire[31:0] T1733;
  wire[31:0] T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire[31:0] T1738;
  wire[31:0] T1739;
  wire[31:0] bankToPort_4_18;
  wire[31:0] T1740;
  wire[31:0] T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire[31:0] T1745;
  wire[31:0] T1746;
  wire[31:0] bankToPort_3_18;
  wire[31:0] T1747;
  wire[31:0] T1748;
  wire T1749;
  wire T1750;
  wire T1751;
  wire[31:0] T1752;
  wire[31:0] T1753;
  wire[31:0] bankToPort_2_18;
  wire[31:0] T1754;
  wire[31:0] T1755;
  wire T1756;
  wire T1757;
  wire T1758;
  wire[31:0] T1759;
  wire[31:0] T1760;
  wire[31:0] bankToPort_1_18;
  wire[31:0] T1761;
  wire[31:0] T1762;
  wire T1763;
  wire T1764;
  wire T1765;
  wire[31:0] T1766;
  wire[31:0] T1767;
  wire[31:0] bankToPort_0_18;
  wire[31:0] T1768;
  wire[31:0] T1769;
  wire T1770;
  wire T1771;
  wire T1772;
  wire T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire[31:0] T1778;
  wire[31:0] T1779;
  wire[31:0] T1780;
  wire[31:0] T1781;
  wire[31:0] T1782;
  wire[31:0] T1783;
  wire[31:0] bankToPort_7_17;
  wire[31:0] T1784;
  wire[31:0] T1785;
  wire T1786;
  wire T1787;
  wire T1788;
  wire[31:0] T1789;
  wire[31:0] T1790;
  wire[31:0] bankToPort_6_17;
  wire[31:0] T1791;
  wire[31:0] T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire[31:0] T1796;
  wire[31:0] T1797;
  wire[31:0] bankToPort_5_17;
  wire[31:0] T1798;
  wire[31:0] T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire[31:0] T1803;
  wire[31:0] T1804;
  wire[31:0] bankToPort_4_17;
  wire[31:0] T1805;
  wire[31:0] T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire[31:0] T1810;
  wire[31:0] T1811;
  wire[31:0] bankToPort_3_17;
  wire[31:0] T1812;
  wire[31:0] T1813;
  wire T1814;
  wire T1815;
  wire T1816;
  wire[31:0] T1817;
  wire[31:0] T1818;
  wire[31:0] bankToPort_2_17;
  wire[31:0] T1819;
  wire[31:0] T1820;
  wire T1821;
  wire T1822;
  wire T1823;
  wire[31:0] T1824;
  wire[31:0] T1825;
  wire[31:0] bankToPort_1_17;
  wire[31:0] T1826;
  wire[31:0] T1827;
  wire T1828;
  wire T1829;
  wire T1830;
  wire[31:0] T1831;
  wire[31:0] T1832;
  wire[31:0] bankToPort_0_17;
  wire[31:0] T1833;
  wire[31:0] T1834;
  wire T1835;
  wire T1836;
  wire T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire T1842;
  wire[31:0] T1843;
  wire[31:0] T1844;
  wire[31:0] T1845;
  wire[31:0] T1846;
  wire[31:0] T1847;
  wire[31:0] T1848;
  wire[31:0] bankToPort_7_16;
  wire[31:0] T1849;
  wire[31:0] T1850;
  wire T1851;
  wire T1852;
  wire T1853;
  wire[31:0] T1854;
  wire[31:0] T1855;
  wire[31:0] bankToPort_6_16;
  wire[31:0] T1856;
  wire[31:0] T1857;
  wire T1858;
  wire T1859;
  wire T1860;
  wire[31:0] T1861;
  wire[31:0] T1862;
  wire[31:0] bankToPort_5_16;
  wire[31:0] T1863;
  wire[31:0] T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[31:0] T1868;
  wire[31:0] T1869;
  wire[31:0] bankToPort_4_16;
  wire[31:0] T1870;
  wire[31:0] T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire[31:0] T1875;
  wire[31:0] T1876;
  wire[31:0] bankToPort_3_16;
  wire[31:0] T1877;
  wire[31:0] T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire[31:0] T1882;
  wire[31:0] T1883;
  wire[31:0] bankToPort_2_16;
  wire[31:0] T1884;
  wire[31:0] T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire[31:0] T1889;
  wire[31:0] T1890;
  wire[31:0] bankToPort_1_16;
  wire[31:0] T1891;
  wire[31:0] T1892;
  wire T1893;
  wire T1894;
  wire T1895;
  wire[31:0] T1896;
  wire[31:0] T1897;
  wire[31:0] bankToPort_0_16;
  wire[31:0] T1898;
  wire[31:0] T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire T1905;
  wire T1906;
  wire T1907;
  wire[31:0] T1908;
  wire[31:0] T1909;
  wire[31:0] T1910;
  wire[31:0] T1911;
  wire[31:0] T1912;
  wire[31:0] T1913;
  wire[31:0] bankToPort_7_15;
  wire[31:0] T1914;
  wire[31:0] T1915;
  wire T1916;
  wire T1917;
  wire T1918;
  wire[31:0] T1919;
  wire[31:0] T1920;
  wire[31:0] bankToPort_6_15;
  wire[31:0] T1921;
  wire[31:0] T1922;
  wire T1923;
  wire T1924;
  wire T1925;
  wire[31:0] T1926;
  wire[31:0] T1927;
  wire[31:0] bankToPort_5_15;
  wire[31:0] T1928;
  wire[31:0] T1929;
  wire T1930;
  wire T1931;
  wire T1932;
  wire[31:0] T1933;
  wire[31:0] T1934;
  wire[31:0] bankToPort_4_15;
  wire[31:0] T1935;
  wire[31:0] T1936;
  wire T1937;
  wire T1938;
  wire T1939;
  wire[31:0] T1940;
  wire[31:0] T1941;
  wire[31:0] bankToPort_3_15;
  wire[31:0] T1942;
  wire[31:0] T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire[31:0] T1947;
  wire[31:0] T1948;
  wire[31:0] bankToPort_2_15;
  wire[31:0] T1949;
  wire[31:0] T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire[31:0] T1954;
  wire[31:0] T1955;
  wire[31:0] bankToPort_1_15;
  wire[31:0] T1956;
  wire[31:0] T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire[31:0] T1961;
  wire[31:0] T1962;
  wire[31:0] bankToPort_0_15;
  wire[31:0] T1963;
  wire[31:0] T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  wire[31:0] T1973;
  wire[31:0] T1974;
  wire[31:0] T1975;
  wire[31:0] T1976;
  wire[31:0] T1977;
  wire[31:0] T1978;
  wire[31:0] bankToPort_7_14;
  wire[31:0] T1979;
  wire[31:0] T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire[31:0] T1984;
  wire[31:0] T1985;
  wire[31:0] bankToPort_6_14;
  wire[31:0] T1986;
  wire[31:0] T1987;
  wire T1988;
  wire T1989;
  wire T1990;
  wire[31:0] T1991;
  wire[31:0] T1992;
  wire[31:0] bankToPort_5_14;
  wire[31:0] T1993;
  wire[31:0] T1994;
  wire T1995;
  wire T1996;
  wire T1997;
  wire[31:0] T1998;
  wire[31:0] T1999;
  wire[31:0] bankToPort_4_14;
  wire[31:0] T2000;
  wire[31:0] T2001;
  wire T2002;
  wire T2003;
  wire T2004;
  wire[31:0] T2005;
  wire[31:0] T2006;
  wire[31:0] bankToPort_3_14;
  wire[31:0] T2007;
  wire[31:0] T2008;
  wire T2009;
  wire T2010;
  wire T2011;
  wire[31:0] T2012;
  wire[31:0] T2013;
  wire[31:0] bankToPort_2_14;
  wire[31:0] T2014;
  wire[31:0] T2015;
  wire T2016;
  wire T2017;
  wire T2018;
  wire[31:0] T2019;
  wire[31:0] T2020;
  wire[31:0] bankToPort_1_14;
  wire[31:0] T2021;
  wire[31:0] T2022;
  wire T2023;
  wire T2024;
  wire T2025;
  wire[31:0] T2026;
  wire[31:0] T2027;
  wire[31:0] bankToPort_0_14;
  wire[31:0] T2028;
  wire[31:0] T2029;
  wire T2030;
  wire T2031;
  wire T2032;
  wire T2033;
  wire T2034;
  wire T2035;
  wire T2036;
  wire T2037;
  wire[31:0] T2038;
  wire[31:0] T2039;
  wire[31:0] T2040;
  wire[31:0] T2041;
  wire[31:0] T2042;
  wire[31:0] T2043;
  wire[31:0] bankToPort_7_13;
  wire[31:0] T2044;
  wire[31:0] T2045;
  wire T2046;
  wire T2047;
  wire T2048;
  wire[31:0] T2049;
  wire[31:0] T2050;
  wire[31:0] bankToPort_6_13;
  wire[31:0] T2051;
  wire[31:0] T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire[31:0] T2056;
  wire[31:0] T2057;
  wire[31:0] bankToPort_5_13;
  wire[31:0] T2058;
  wire[31:0] T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire[31:0] T2063;
  wire[31:0] T2064;
  wire[31:0] bankToPort_4_13;
  wire[31:0] T2065;
  wire[31:0] T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire[31:0] T2070;
  wire[31:0] T2071;
  wire[31:0] bankToPort_3_13;
  wire[31:0] T2072;
  wire[31:0] T2073;
  wire T2074;
  wire T2075;
  wire T2076;
  wire[31:0] T2077;
  wire[31:0] T2078;
  wire[31:0] bankToPort_2_13;
  wire[31:0] T2079;
  wire[31:0] T2080;
  wire T2081;
  wire T2082;
  wire T2083;
  wire[31:0] T2084;
  wire[31:0] T2085;
  wire[31:0] bankToPort_1_13;
  wire[31:0] T2086;
  wire[31:0] T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire[31:0] T2091;
  wire[31:0] T2092;
  wire[31:0] bankToPort_0_13;
  wire[31:0] T2093;
  wire[31:0] T2094;
  wire T2095;
  wire T2096;
  wire T2097;
  wire T2098;
  wire T2099;
  wire T2100;
  wire T2101;
  wire T2102;
  wire[31:0] T2103;
  wire[31:0] T2104;
  wire[31:0] T2105;
  wire[31:0] T2106;
  wire[31:0] T2107;
  wire[31:0] T2108;
  wire[31:0] bankToPort_7_12;
  wire[31:0] T2109;
  wire[31:0] T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire[31:0] T2114;
  wire[31:0] T2115;
  wire[31:0] bankToPort_6_12;
  wire[31:0] T2116;
  wire[31:0] T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[31:0] T2121;
  wire[31:0] T2122;
  wire[31:0] bankToPort_5_12;
  wire[31:0] T2123;
  wire[31:0] T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire[31:0] T2128;
  wire[31:0] T2129;
  wire[31:0] bankToPort_4_12;
  wire[31:0] T2130;
  wire[31:0] T2131;
  wire T2132;
  wire T2133;
  wire T2134;
  wire[31:0] T2135;
  wire[31:0] T2136;
  wire[31:0] bankToPort_3_12;
  wire[31:0] T2137;
  wire[31:0] T2138;
  wire T2139;
  wire T2140;
  wire T2141;
  wire[31:0] T2142;
  wire[31:0] T2143;
  wire[31:0] bankToPort_2_12;
  wire[31:0] T2144;
  wire[31:0] T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire[31:0] T2149;
  wire[31:0] T2150;
  wire[31:0] bankToPort_1_12;
  wire[31:0] T2151;
  wire[31:0] T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire[31:0] T2156;
  wire[31:0] T2157;
  wire[31:0] bankToPort_0_12;
  wire[31:0] T2158;
  wire[31:0] T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  wire T2165;
  wire T2166;
  wire T2167;
  wire[31:0] T2168;
  wire[31:0] T2169;
  wire[31:0] T2170;
  wire[31:0] T2171;
  wire[31:0] T2172;
  wire[31:0] T2173;
  wire[31:0] bankToPort_7_11;
  wire[31:0] T2174;
  wire[31:0] T2175;
  wire T2176;
  wire T2177;
  wire T2178;
  wire[31:0] T2179;
  wire[31:0] T2180;
  wire[31:0] bankToPort_6_11;
  wire[31:0] T2181;
  wire[31:0] T2182;
  wire T2183;
  wire T2184;
  wire T2185;
  wire[31:0] T2186;
  wire[31:0] T2187;
  wire[31:0] bankToPort_5_11;
  wire[31:0] T2188;
  wire[31:0] T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[31:0] T2193;
  wire[31:0] T2194;
  wire[31:0] bankToPort_4_11;
  wire[31:0] T2195;
  wire[31:0] T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire[31:0] T2200;
  wire[31:0] T2201;
  wire[31:0] bankToPort_3_11;
  wire[31:0] T2202;
  wire[31:0] T2203;
  wire T2204;
  wire T2205;
  wire T2206;
  wire[31:0] T2207;
  wire[31:0] T2208;
  wire[31:0] bankToPort_2_11;
  wire[31:0] T2209;
  wire[31:0] T2210;
  wire T2211;
  wire T2212;
  wire T2213;
  wire[31:0] T2214;
  wire[31:0] T2215;
  wire[31:0] bankToPort_1_11;
  wire[31:0] T2216;
  wire[31:0] T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  wire[31:0] T2221;
  wire[31:0] T2222;
  wire[31:0] bankToPort_0_11;
  wire[31:0] T2223;
  wire[31:0] T2224;
  wire T2225;
  wire T2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire[31:0] T2233;
  wire[31:0] T2234;
  wire[31:0] T2235;
  wire[31:0] T2236;
  wire[31:0] T2237;
  wire[31:0] T2238;
  wire[31:0] bankToPort_7_10;
  wire[31:0] T2239;
  wire[31:0] T2240;
  wire T2241;
  wire T2242;
  wire T2243;
  wire[31:0] T2244;
  wire[31:0] T2245;
  wire[31:0] bankToPort_6_10;
  wire[31:0] T2246;
  wire[31:0] T2247;
  wire T2248;
  wire T2249;
  wire T2250;
  wire[31:0] T2251;
  wire[31:0] T2252;
  wire[31:0] bankToPort_5_10;
  wire[31:0] T2253;
  wire[31:0] T2254;
  wire T2255;
  wire T2256;
  wire T2257;
  wire[31:0] T2258;
  wire[31:0] T2259;
  wire[31:0] bankToPort_4_10;
  wire[31:0] T2260;
  wire[31:0] T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[31:0] T2265;
  wire[31:0] T2266;
  wire[31:0] bankToPort_3_10;
  wire[31:0] T2267;
  wire[31:0] T2268;
  wire T2269;
  wire T2270;
  wire T2271;
  wire[31:0] T2272;
  wire[31:0] T2273;
  wire[31:0] bankToPort_2_10;
  wire[31:0] T2274;
  wire[31:0] T2275;
  wire T2276;
  wire T2277;
  wire T2278;
  wire[31:0] T2279;
  wire[31:0] T2280;
  wire[31:0] bankToPort_1_10;
  wire[31:0] T2281;
  wire[31:0] T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  wire[31:0] T2286;
  wire[31:0] T2287;
  wire[31:0] bankToPort_0_10;
  wire[31:0] T2288;
  wire[31:0] T2289;
  wire T2290;
  wire T2291;
  wire T2292;
  wire T2293;
  wire T2294;
  wire T2295;
  wire T2296;
  wire T2297;
  wire[31:0] T2298;
  wire[31:0] T2299;
  wire[31:0] T2300;
  wire[31:0] T2301;
  wire[31:0] T2302;
  wire[31:0] T2303;
  wire[31:0] bankToPort_7_9;
  wire[31:0] T2304;
  wire[31:0] T2305;
  wire T2306;
  wire T2307;
  wire T2308;
  wire[31:0] T2309;
  wire[31:0] T2310;
  wire[31:0] bankToPort_6_9;
  wire[31:0] T2311;
  wire[31:0] T2312;
  wire T2313;
  wire T2314;
  wire T2315;
  wire[31:0] T2316;
  wire[31:0] T2317;
  wire[31:0] bankToPort_5_9;
  wire[31:0] T2318;
  wire[31:0] T2319;
  wire T2320;
  wire T2321;
  wire T2322;
  wire[31:0] T2323;
  wire[31:0] T2324;
  wire[31:0] bankToPort_4_9;
  wire[31:0] T2325;
  wire[31:0] T2326;
  wire T2327;
  wire T2328;
  wire T2329;
  wire[31:0] T2330;
  wire[31:0] T2331;
  wire[31:0] bankToPort_3_9;
  wire[31:0] T2332;
  wire[31:0] T2333;
  wire T2334;
  wire T2335;
  wire T2336;
  wire[31:0] T2337;
  wire[31:0] T2338;
  wire[31:0] bankToPort_2_9;
  wire[31:0] T2339;
  wire[31:0] T2340;
  wire T2341;
  wire T2342;
  wire T2343;
  wire[31:0] T2344;
  wire[31:0] T2345;
  wire[31:0] bankToPort_1_9;
  wire[31:0] T2346;
  wire[31:0] T2347;
  wire T2348;
  wire T2349;
  wire T2350;
  wire[31:0] T2351;
  wire[31:0] T2352;
  wire[31:0] bankToPort_0_9;
  wire[31:0] T2353;
  wire[31:0] T2354;
  wire T2355;
  wire T2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  wire T2361;
  wire T2362;
  wire[31:0] T2363;
  wire[31:0] T2364;
  wire[31:0] T2365;
  wire[31:0] T2366;
  wire[31:0] T2367;
  wire[31:0] T2368;
  wire[31:0] bankToPort_7_8;
  wire[31:0] T2369;
  wire[31:0] T2370;
  wire T2371;
  wire T2372;
  wire T2373;
  wire[31:0] T2374;
  wire[31:0] T2375;
  wire[31:0] bankToPort_6_8;
  wire[31:0] T2376;
  wire[31:0] T2377;
  wire T2378;
  wire T2379;
  wire T2380;
  wire[31:0] T2381;
  wire[31:0] T2382;
  wire[31:0] bankToPort_5_8;
  wire[31:0] T2383;
  wire[31:0] T2384;
  wire T2385;
  wire T2386;
  wire T2387;
  wire[31:0] T2388;
  wire[31:0] T2389;
  wire[31:0] bankToPort_4_8;
  wire[31:0] T2390;
  wire[31:0] T2391;
  wire T2392;
  wire T2393;
  wire T2394;
  wire[31:0] T2395;
  wire[31:0] T2396;
  wire[31:0] bankToPort_3_8;
  wire[31:0] T2397;
  wire[31:0] T2398;
  wire T2399;
  wire T2400;
  wire T2401;
  wire[31:0] T2402;
  wire[31:0] T2403;
  wire[31:0] bankToPort_2_8;
  wire[31:0] T2404;
  wire[31:0] T2405;
  wire T2406;
  wire T2407;
  wire T2408;
  wire[31:0] T2409;
  wire[31:0] T2410;
  wire[31:0] bankToPort_1_8;
  wire[31:0] T2411;
  wire[31:0] T2412;
  wire T2413;
  wire T2414;
  wire T2415;
  wire[31:0] T2416;
  wire[31:0] T2417;
  wire[31:0] bankToPort_0_8;
  wire[31:0] T2418;
  wire[31:0] T2419;
  wire T2420;
  wire T2421;
  wire T2422;
  wire T2423;
  wire T2424;
  wire T2425;
  wire T2426;
  wire T2427;
  wire[31:0] T2428;
  wire[31:0] T2429;
  wire[31:0] T2430;
  wire[31:0] T2431;
  wire[31:0] T2432;
  wire[31:0] T2433;
  wire[31:0] bankToPort_7_7;
  wire[31:0] T2434;
  wire[31:0] T2435;
  wire T2436;
  wire T2437;
  wire T2438;
  wire[31:0] T2439;
  wire[31:0] T2440;
  wire[31:0] bankToPort_6_7;
  wire[31:0] T2441;
  wire[31:0] T2442;
  wire T2443;
  wire T2444;
  wire T2445;
  wire[31:0] T2446;
  wire[31:0] T2447;
  wire[31:0] bankToPort_5_7;
  wire[31:0] T2448;
  wire[31:0] T2449;
  wire T2450;
  wire T2451;
  wire T2452;
  wire[31:0] T2453;
  wire[31:0] T2454;
  wire[31:0] bankToPort_4_7;
  wire[31:0] T2455;
  wire[31:0] T2456;
  wire T2457;
  wire T2458;
  wire T2459;
  wire[31:0] T2460;
  wire[31:0] T2461;
  wire[31:0] bankToPort_3_7;
  wire[31:0] T2462;
  wire[31:0] T2463;
  wire T2464;
  wire T2465;
  wire T2466;
  wire[31:0] T2467;
  wire[31:0] T2468;
  wire[31:0] bankToPort_2_7;
  wire[31:0] T2469;
  wire[31:0] T2470;
  wire T2471;
  wire T2472;
  wire T2473;
  wire[31:0] T2474;
  wire[31:0] T2475;
  wire[31:0] bankToPort_1_7;
  wire[31:0] T2476;
  wire[31:0] T2477;
  wire T2478;
  wire T2479;
  wire T2480;
  wire[31:0] T2481;
  wire[31:0] T2482;
  wire[31:0] bankToPort_0_7;
  wire[31:0] T2483;
  wire[31:0] T2484;
  wire T2485;
  wire T2486;
  wire T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  wire T2491;
  wire T2492;
  wire[31:0] T2493;
  wire[31:0] T2494;
  wire[31:0] T2495;
  wire[31:0] T2496;
  wire[31:0] T2497;
  wire[31:0] T2498;
  wire[31:0] bankToPort_7_6;
  wire[31:0] T2499;
  wire[31:0] T2500;
  wire T2501;
  wire T2502;
  wire T2503;
  wire[31:0] T2504;
  wire[31:0] T2505;
  wire[31:0] bankToPort_6_6;
  wire[31:0] T2506;
  wire[31:0] T2507;
  wire T2508;
  wire T2509;
  wire T2510;
  wire[31:0] T2511;
  wire[31:0] T2512;
  wire[31:0] bankToPort_5_6;
  wire[31:0] T2513;
  wire[31:0] T2514;
  wire T2515;
  wire T2516;
  wire T2517;
  wire[31:0] T2518;
  wire[31:0] T2519;
  wire[31:0] bankToPort_4_6;
  wire[31:0] T2520;
  wire[31:0] T2521;
  wire T2522;
  wire T2523;
  wire T2524;
  wire[31:0] T2525;
  wire[31:0] T2526;
  wire[31:0] bankToPort_3_6;
  wire[31:0] T2527;
  wire[31:0] T2528;
  wire T2529;
  wire T2530;
  wire T2531;
  wire[31:0] T2532;
  wire[31:0] T2533;
  wire[31:0] bankToPort_2_6;
  wire[31:0] T2534;
  wire[31:0] T2535;
  wire T2536;
  wire T2537;
  wire T2538;
  wire[31:0] T2539;
  wire[31:0] T2540;
  wire[31:0] bankToPort_1_6;
  wire[31:0] T2541;
  wire[31:0] T2542;
  wire T2543;
  wire T2544;
  wire T2545;
  wire[31:0] T2546;
  wire[31:0] T2547;
  wire[31:0] bankToPort_0_6;
  wire[31:0] T2548;
  wire[31:0] T2549;
  wire T2550;
  wire T2551;
  wire T2552;
  wire T2553;
  wire T2554;
  wire T2555;
  wire T2556;
  wire T2557;
  wire[31:0] T2558;
  wire[31:0] T2559;
  wire[31:0] T2560;
  wire[31:0] T2561;
  wire[31:0] T2562;
  wire[31:0] T2563;
  wire[31:0] bankToPort_7_5;
  wire[31:0] T2564;
  wire[31:0] T2565;
  wire T2566;
  wire T2567;
  wire T2568;
  wire[31:0] T2569;
  wire[31:0] T2570;
  wire[31:0] bankToPort_6_5;
  wire[31:0] T2571;
  wire[31:0] T2572;
  wire T2573;
  wire T2574;
  wire T2575;
  wire[31:0] T2576;
  wire[31:0] T2577;
  wire[31:0] bankToPort_5_5;
  wire[31:0] T2578;
  wire[31:0] T2579;
  wire T2580;
  wire T2581;
  wire T2582;
  wire[31:0] T2583;
  wire[31:0] T2584;
  wire[31:0] bankToPort_4_5;
  wire[31:0] T2585;
  wire[31:0] T2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire[31:0] T2590;
  wire[31:0] T2591;
  wire[31:0] bankToPort_3_5;
  wire[31:0] T2592;
  wire[31:0] T2593;
  wire T2594;
  wire T2595;
  wire T2596;
  wire[31:0] T2597;
  wire[31:0] T2598;
  wire[31:0] bankToPort_2_5;
  wire[31:0] T2599;
  wire[31:0] T2600;
  wire T2601;
  wire T2602;
  wire T2603;
  wire[31:0] T2604;
  wire[31:0] T2605;
  wire[31:0] bankToPort_1_5;
  wire[31:0] T2606;
  wire[31:0] T2607;
  wire T2608;
  wire T2609;
  wire T2610;
  wire[31:0] T2611;
  wire[31:0] T2612;
  wire[31:0] bankToPort_0_5;
  wire[31:0] T2613;
  wire[31:0] T2614;
  wire T2615;
  wire T2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire T2620;
  wire T2621;
  wire T2622;
  wire[31:0] T2623;
  wire[31:0] T2624;
  wire[31:0] T2625;
  wire[31:0] T2626;
  wire[31:0] T2627;
  wire[31:0] T2628;
  wire[31:0] bankToPort_7_4;
  wire[31:0] T2629;
  wire[31:0] T2630;
  wire T2631;
  wire T2632;
  wire T2633;
  wire[31:0] T2634;
  wire[31:0] T2635;
  wire[31:0] bankToPort_6_4;
  wire[31:0] T2636;
  wire[31:0] T2637;
  wire T2638;
  wire T2639;
  wire T2640;
  wire[31:0] T2641;
  wire[31:0] T2642;
  wire[31:0] bankToPort_5_4;
  wire[31:0] T2643;
  wire[31:0] T2644;
  wire T2645;
  wire T2646;
  wire T2647;
  wire[31:0] T2648;
  wire[31:0] T2649;
  wire[31:0] bankToPort_4_4;
  wire[31:0] T2650;
  wire[31:0] T2651;
  wire T2652;
  wire T2653;
  wire T2654;
  wire[31:0] T2655;
  wire[31:0] T2656;
  wire[31:0] bankToPort_3_4;
  wire[31:0] T2657;
  wire[31:0] T2658;
  wire T2659;
  wire T2660;
  wire T2661;
  wire[31:0] T2662;
  wire[31:0] T2663;
  wire[31:0] bankToPort_2_4;
  wire[31:0] T2664;
  wire[31:0] T2665;
  wire T2666;
  wire T2667;
  wire T2668;
  wire[31:0] T2669;
  wire[31:0] T2670;
  wire[31:0] bankToPort_1_4;
  wire[31:0] T2671;
  wire[31:0] T2672;
  wire T2673;
  wire T2674;
  wire T2675;
  wire[31:0] T2676;
  wire[31:0] T2677;
  wire[31:0] bankToPort_0_4;
  wire[31:0] T2678;
  wire[31:0] T2679;
  wire T2680;
  wire T2681;
  wire T2682;
  wire T2683;
  wire T2684;
  wire T2685;
  wire T2686;
  wire T2687;
  wire[31:0] T2688;
  wire[31:0] T2689;
  wire[31:0] T2690;
  wire[31:0] T2691;
  wire[31:0] T2692;
  wire[31:0] T2693;
  wire[31:0] bankToPort_7_3;
  wire[31:0] T2694;
  wire[31:0] T2695;
  wire T2696;
  wire T2697;
  wire T2698;
  wire[31:0] T2699;
  wire[31:0] T2700;
  wire[31:0] bankToPort_6_3;
  wire[31:0] T2701;
  wire[31:0] T2702;
  wire T2703;
  wire T2704;
  wire T2705;
  wire[31:0] T2706;
  wire[31:0] T2707;
  wire[31:0] bankToPort_5_3;
  wire[31:0] T2708;
  wire[31:0] T2709;
  wire T2710;
  wire T2711;
  wire T2712;
  wire[31:0] T2713;
  wire[31:0] T2714;
  wire[31:0] bankToPort_4_3;
  wire[31:0] T2715;
  wire[31:0] T2716;
  wire T2717;
  wire T2718;
  wire T2719;
  wire[31:0] T2720;
  wire[31:0] T2721;
  wire[31:0] bankToPort_3_3;
  wire[31:0] T2722;
  wire[31:0] T2723;
  wire T2724;
  wire T2725;
  wire T2726;
  wire[31:0] T2727;
  wire[31:0] T2728;
  wire[31:0] bankToPort_2_3;
  wire[31:0] T2729;
  wire[31:0] T2730;
  wire T2731;
  wire T2732;
  wire T2733;
  wire[31:0] T2734;
  wire[31:0] T2735;
  wire[31:0] bankToPort_1_3;
  wire[31:0] T2736;
  wire[31:0] T2737;
  wire T2738;
  wire T2739;
  wire T2740;
  wire[31:0] T2741;
  wire[31:0] T2742;
  wire[31:0] bankToPort_0_3;
  wire[31:0] T2743;
  wire[31:0] T2744;
  wire T2745;
  wire T2746;
  wire T2747;
  wire T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  wire T2752;
  wire[31:0] T2753;
  wire[31:0] T2754;
  wire[31:0] T2755;
  wire[31:0] T2756;
  wire[31:0] T2757;
  wire[31:0] T2758;
  wire[31:0] bankToPort_7_2;
  wire[31:0] T2759;
  wire[31:0] T2760;
  wire T2761;
  wire T2762;
  wire T2763;
  wire[31:0] T2764;
  wire[31:0] T2765;
  wire[31:0] bankToPort_6_2;
  wire[31:0] T2766;
  wire[31:0] T2767;
  wire T2768;
  wire T2769;
  wire T2770;
  wire[31:0] T2771;
  wire[31:0] T2772;
  wire[31:0] bankToPort_5_2;
  wire[31:0] T2773;
  wire[31:0] T2774;
  wire T2775;
  wire T2776;
  wire T2777;
  wire[31:0] T2778;
  wire[31:0] T2779;
  wire[31:0] bankToPort_4_2;
  wire[31:0] T2780;
  wire[31:0] T2781;
  wire T2782;
  wire T2783;
  wire T2784;
  wire[31:0] T2785;
  wire[31:0] T2786;
  wire[31:0] bankToPort_3_2;
  wire[31:0] T2787;
  wire[31:0] T2788;
  wire T2789;
  wire T2790;
  wire T2791;
  wire[31:0] T2792;
  wire[31:0] T2793;
  wire[31:0] bankToPort_2_2;
  wire[31:0] T2794;
  wire[31:0] T2795;
  wire T2796;
  wire T2797;
  wire T2798;
  wire[31:0] T2799;
  wire[31:0] T2800;
  wire[31:0] bankToPort_1_2;
  wire[31:0] T2801;
  wire[31:0] T2802;
  wire T2803;
  wire T2804;
  wire T2805;
  wire[31:0] T2806;
  wire[31:0] T2807;
  wire[31:0] bankToPort_0_2;
  wire[31:0] T2808;
  wire[31:0] T2809;
  wire T2810;
  wire T2811;
  wire T2812;
  wire T2813;
  wire T2814;
  wire T2815;
  wire T2816;
  wire T2817;
  wire[31:0] T2818;
  wire[31:0] T2819;
  wire[31:0] T2820;
  wire[31:0] T2821;
  wire[31:0] T2822;
  wire[31:0] T2823;
  wire[31:0] bankToPort_7_1;
  wire[31:0] T2824;
  wire[31:0] T2825;
  wire T2826;
  wire T2827;
  wire T2828;
  wire[31:0] T2829;
  wire[31:0] T2830;
  wire[31:0] bankToPort_6_1;
  wire[31:0] T2831;
  wire[31:0] T2832;
  wire T2833;
  wire T2834;
  wire T2835;
  wire[31:0] T2836;
  wire[31:0] T2837;
  wire[31:0] bankToPort_5_1;
  wire[31:0] T2838;
  wire[31:0] T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  wire[31:0] T2843;
  wire[31:0] T2844;
  wire[31:0] bankToPort_4_1;
  wire[31:0] T2845;
  wire[31:0] T2846;
  wire T2847;
  wire T2848;
  wire T2849;
  wire[31:0] T2850;
  wire[31:0] T2851;
  wire[31:0] bankToPort_3_1;
  wire[31:0] T2852;
  wire[31:0] T2853;
  wire T2854;
  wire T2855;
  wire T2856;
  wire[31:0] T2857;
  wire[31:0] T2858;
  wire[31:0] bankToPort_2_1;
  wire[31:0] T2859;
  wire[31:0] T2860;
  wire T2861;
  wire T2862;
  wire T2863;
  wire[31:0] T2864;
  wire[31:0] T2865;
  wire[31:0] bankToPort_1_1;
  wire[31:0] T2866;
  wire[31:0] T2867;
  wire T2868;
  wire T2869;
  wire T2870;
  wire[31:0] T2871;
  wire[31:0] T2872;
  wire[31:0] bankToPort_0_1;
  wire[31:0] T2873;
  wire[31:0] T2874;
  wire T2875;
  wire T2876;
  wire T2877;
  wire T2878;
  wire T2879;
  wire T2880;
  wire T2881;
  wire T2882;
  wire[31:0] T2883;
  wire[31:0] T2884;
  wire[31:0] T2885;
  wire[31:0] T2886;
  wire[31:0] T2887;
  wire[31:0] T2888;
  wire[31:0] bankToPort_7_0;
  wire[31:0] T2889;
  wire[31:0] T2890;
  wire T2891;
  wire T2892;
  wire T2893;
  wire[31:0] T2894;
  wire[31:0] T2895;
  wire[31:0] bankToPort_6_0;
  wire[31:0] T2896;
  wire[31:0] T2897;
  wire T2898;
  wire T2899;
  wire T2900;
  wire[31:0] T2901;
  wire[31:0] T2902;
  wire[31:0] bankToPort_5_0;
  wire[31:0] T2903;
  wire[31:0] T2904;
  wire T2905;
  wire T2906;
  wire T2907;
  wire[31:0] T2908;
  wire[31:0] T2909;
  wire[31:0] bankToPort_4_0;
  wire[31:0] T2910;
  wire[31:0] T2911;
  wire T2912;
  wire T2913;
  wire T2914;
  wire[31:0] T2915;
  wire[31:0] T2916;
  wire[31:0] bankToPort_3_0;
  wire[31:0] T2917;
  wire[31:0] T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire[31:0] T2922;
  wire[31:0] T2923;
  wire[31:0] bankToPort_2_0;
  wire[31:0] T2924;
  wire[31:0] T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire[31:0] T2929;
  wire[31:0] T2930;
  wire[31:0] bankToPort_1_0;
  wire[31:0] T2931;
  wire[31:0] T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire[31:0] T2936;
  wire[31:0] T2937;
  wire[31:0] bankToPort_0_0;
  wire[31:0] T2938;
  wire[31:0] T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire T2943;
  wire T2944;
  wire T2945;
  wire[31:0] T2946;
  wire T2947;
  wire T2948;
  wire[31:0] T2949;
  wire T2950;
  wire T2951;
  wire[31:0] T2952;
  wire T2953;
  wire T2954;
  wire[31:0] T2955;
  wire T2956;
  wire T2957;
  wire[31:0] T2958;
  wire T2959;
  wire T2960;
  wire[31:0] T2961;
  wire T2962;
  wire T2963;
  wire[31:0] T2964;
  wire T2965;
  wire T2966;
  wire[31:0] T2967;
  wire T2968;
  wire T2969;
  wire[31:0] T2970;
  wire T2971;
  wire T2972;
  wire[31:0] T2973;
  wire T2974;
  wire T2975;
  wire[31:0] T2976;
  wire T2977;
  wire T2978;
  wire[31:0] T2979;
  wire T2980;
  wire T2981;
  wire[31:0] T2982;
  wire T2983;
  wire T2984;
  wire[31:0] T2985;
  wire T2986;
  wire T2987;
  wire[31:0] T2988;
  wire T2989;
  wire T2990;
  wire[31:0] T2991;
  wire T2992;
  wire T2993;
  wire[31:0] T2994;
  wire T2995;
  wire T2996;
  wire[31:0] T2997;
  wire T2998;
  wire T2999;
  wire[31:0] T3000;
  wire T3001;
  wire T3002;
  wire[31:0] T3003;
  wire T3004;
  wire T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire T3013;
  wire T3014;
  wire T3015;
  wire T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire T3028;
  wire T3029;
  wire T3030;
  wire T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire T3043;
  wire T3044;
  wire T3045;
  wire T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire T3050;
  wire T3051;
  wire T3052;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire T3057;
  wire T3058;
  wire T3059;
  wire T3060;
  wire[5:0] T3061;
  wire[5:0] readAddr;
  wire[5:0] T3062;
  wire[5:0] T3063;
  wire[5:0] T3064;
  wire[5:0] T3065;
  wire[5:0] T3066;
  wire[5:0] T3067;
  wire[5:0] T3068;
  wire[5:0] T3069;
  wire[5:0] T3070;
  wire[5:0] T3071;
  wire[5:0] T3072;
  wire[5:0] T3073;
  wire[5:0] T3074;
  wire[5:0] T3075;
  wire[5:0] T3076;
  wire[5:0] T3077;
  wire[5:0] T3078;
  wire[5:0] T3079;
  wire[5:0] T3080;
  wire[5:0] T3081;
  wire[5:0] T3082;
  wire[5:0] T3083;
  wire[5:0] T3084;
  wire[5:0] T3085;
  wire[5:0] T3086;
  wire[5:0] T3087;
  wire[5:0] T3088;
  wire[5:0] T3089;
  wire[5:0] T3090;
  wire[5:0] T3091;
  wire[8:0] T3092;
  wire T3093;
  wire T3094;
  wire T3095;
  wire T3096;
  wire T3097;
  wire[88:0] fabInSeqMem_io_outData;
  wire[8:0] fabInSeqMemConfig_io_memAddr;
  wire[88:0] fabInSeqMemConfig_io_memData;
  wire fabInSeqMemConfig_io_memOutValid;
  wire fabInSeqMemConfig_io_rst;
  wire[31:0] fifo_io_deqData;
  wire fifo_io_enqRdy;
  wire fifo_io_deqValid;
  wire[31:0] fifo_1_io_deqData;
  wire fifo_1_io_enqRdy;
  wire fifo_1_io_deqValid;
  wire[31:0] fifo_2_io_deqData;
  wire fifo_2_io_enqRdy;
  wire fifo_2_io_deqValid;
  wire[31:0] fifo_3_io_deqData;
  wire fifo_3_io_enqRdy;
  wire fifo_3_io_deqValid;
  wire[31:0] fifo_4_io_deqData;
  wire fifo_4_io_enqRdy;
  wire fifo_4_io_deqValid;
  wire[31:0] fifo_5_io_deqData;
  wire fifo_5_io_enqRdy;
  wire fifo_5_io_deqValid;
  wire[31:0] fifo_6_io_deqData;
  wire fifo_6_io_enqRdy;
  wire fifo_6_io_deqValid;
  wire[31:0] fifo_7_io_deqData;
  wire fifo_7_io_enqRdy;
  wire fifo_7_io_deqValid;
  wire[31:0] fifo_8_io_deqData;
  wire fifo_8_io_enqRdy;
  wire fifo_8_io_deqValid;
  wire[31:0] fifo_9_io_deqData;
  wire fifo_9_io_enqRdy;
  wire fifo_9_io_deqValid;
  wire[31:0] fifo_10_io_deqData;
  wire fifo_10_io_enqRdy;
  wire fifo_10_io_deqValid;
  wire[31:0] fifo_11_io_deqData;
  wire fifo_11_io_enqRdy;
  wire fifo_11_io_deqValid;
  wire[31:0] fifo_12_io_deqData;
  wire fifo_12_io_enqRdy;
  wire fifo_12_io_deqValid;
  wire[31:0] fifo_13_io_deqData;
  wire fifo_13_io_enqRdy;
  wire fifo_13_io_deqValid;
  wire[31:0] fifo_14_io_deqData;
  wire fifo_14_io_enqRdy;
  wire fifo_14_io_deqValid;
  wire[31:0] fifo_15_io_deqData;
  wire fifo_15_io_enqRdy;
  wire fifo_15_io_deqValid;
  wire[31:0] fifo_16_io_deqData;
  wire fifo_16_io_enqRdy;
  wire fifo_16_io_deqValid;
  wire[31:0] fifo_17_io_deqData;
  wire fifo_17_io_enqRdy;
  wire fifo_17_io_deqValid;
  wire[31:0] fifo_18_io_deqData;
  wire fifo_18_io_enqRdy;
  wire fifo_18_io_deqValid;
  wire[31:0] fifo_19_io_deqData;
  wire fifo_19_io_enqRdy;
  wire fifo_19_io_deqValid;
  wire[31:0] fifo_20_io_deqData;
  wire fifo_20_io_enqRdy;
  wire fifo_20_io_deqValid;
  wire[31:0] fifo_21_io_deqData;
  wire fifo_21_io_enqRdy;
  wire fifo_21_io_deqValid;
  wire[31:0] fifo_22_io_deqData;
  wire fifo_22_io_enqRdy;
  wire fifo_22_io_deqValid;
  wire[31:0] fifo_23_io_deqData;
  wire fifo_23_io_enqRdy;
  wire fifo_23_io_deqValid;
  wire[31:0] fifo_24_io_deqData;
  wire fifo_24_io_enqRdy;
  wire fifo_24_io_deqValid;
  wire[31:0] fifo_25_io_deqData;
  wire fifo_25_io_enqRdy;
  wire fifo_25_io_deqValid;
  wire[31:0] fifo_26_io_deqData;
  wire fifo_26_io_enqRdy;
  wire fifo_26_io_deqValid;
  wire[31:0] fifo_27_io_deqData;
  wire fifo_27_io_enqRdy;
  wire fifo_27_io_deqValid;
  wire[31:0] fifo_28_io_deqData;
  wire fifo_28_io_enqRdy;
  wire fifo_28_io_deqValid;
  wire[31:0] fifo_29_io_deqData;
  wire fifo_29_io_enqRdy;
  wire fifo_29_io_deqValid;
  wire[31:0] fifo_30_io_deqData;
  wire fifo_30_io_enqRdy;
  wire fifo_30_io_deqValid;
  wire[31:0] fifo_31_io_deqData;
  wire fifo_31_io_enqRdy;
  wire fifo_31_io_deqValid;
  wire[31:0] fifo_32_io_deqData;
  wire fifo_32_io_enqRdy;
  wire fifo_32_io_deqValid;
  wire[31:0] fifo_33_io_deqData;
  wire fifo_33_io_enqRdy;
  wire fifo_33_io_deqValid;
  wire[31:0] fifo_34_io_deqData;
  wire fifo_34_io_enqRdy;
  wire fifo_34_io_deqValid;
  wire[31:0] fifo_35_io_deqData;
  wire fifo_35_io_enqRdy;
  wire fifo_35_io_deqValid;
  wire[31:0] fifo_36_io_deqData;
  wire fifo_36_io_enqRdy;
  wire fifo_36_io_deqValid;
  wire[31:0] fifo_37_io_deqData;
  wire fifo_37_io_enqRdy;
  wire fifo_37_io_deqValid;
  wire[31:0] fifo_38_io_deqData;
  wire fifo_38_io_enqRdy;
  wire fifo_38_io_deqValid;
  wire[31:0] fifo_39_io_deqData;
  wire fifo_39_io_enqRdy;
  wire fifo_39_io_deqValid;
  wire[31:0] fifo_40_io_deqData;
  wire fifo_40_io_enqRdy;
  wire fifo_40_io_deqValid;
  wire[31:0] fifo_41_io_deqData;
  wire fifo_41_io_enqRdy;
  wire fifo_41_io_deqValid;
  wire[31:0] fifo_42_io_deqData;
  wire fifo_42_io_enqRdy;
  wire fifo_42_io_deqValid;
  wire[31:0] fifo_43_io_deqData;
  wire fifo_43_io_enqRdy;
  wire fifo_43_io_deqValid;
  wire[31:0] fifo_44_io_deqData;
  wire fifo_44_io_enqRdy;
  wire fifo_44_io_deqValid;
  wire[31:0] fifo_45_io_deqData;
  wire fifo_45_io_enqRdy;
  wire fifo_45_io_deqValid;
  wire[31:0] fifo_46_io_deqData;
  wire fifo_46_io_enqRdy;
  wire fifo_46_io_deqValid;
  wire[31:0] fifo_47_io_deqData;
  wire fifo_47_io_enqRdy;
  wire fifo_47_io_deqValid;
  wire[37:0] localStorage_io_outData_7;
  wire[37:0] localStorage_io_outData_6;
  wire[37:0] localStorage_io_outData_5;
  wire[37:0] localStorage_io_outData_4;
  wire[37:0] localStorage_io_outData_3;
  wire[37:0] localStorage_io_outData_2;
  wire[37:0] localStorage_io_outData_1;
  wire[37:0] localStorage_io_outData_0;
  wire localStorage_io_isReadValid_7;
  wire localStorage_io_isReadValid_6;
  wire localStorage_io_isReadValid_5;
  wire localStorage_io_isReadValid_4;
  wire localStorage_io_isReadValid_3;
  wire localStorage_io_isReadValid_2;
  wire localStorage_io_isReadValid_1;
  wire localStorage_io_isReadValid_0;
  wire localStorage_io_enqRdyLoad_7;
  wire localStorage_io_enqRdyLoad_6;
  wire localStorage_io_enqRdyLoad_5;
  wire localStorage_io_enqRdyLoad_4;
  wire localStorage_io_enqRdyLoad_3;
  wire localStorage_io_enqRdyLoad_2;
  wire localStorage_io_enqRdyLoad_1;
  wire localStorage_io_enqRdyLoad_0;
  wire localStorage_io_enqRdyFabric_7;
  wire localStorage_io_enqRdyFabric_6;
  wire localStorage_io_enqRdyFabric_5;
  wire localStorage_io_enqRdyFabric_4;
  wire localStorage_io_enqRdyFabric_3;
  wire localStorage_io_enqRdyFabric_2;
  wire localStorage_io_enqRdyFabric_1;
  wire localStorage_io_enqRdyFabric_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    nextSeqSelReg = {1{$random}};
    nextSeqReg2 = {3{$random}};
    firstSeqSelReg = {1{$random}};
    bankReadDoneReg_1 = {1{$random}};
    nextSeqRegValid2 = {1{$random}};
    nextSeqRegValid1 = {1{$random}};
    bankReadDoneReg_2 = {1{$random}};
    bankReadDoneReg_3 = {1{$random}};
    bankReadDoneReg_4 = {1{$random}};
    bankReadDoneReg_5 = {1{$random}};
    bankReadDoneReg_6 = {1{$random}};
    bankReadDoneReg_7 = {1{$random}};
    bankReadDoneReg_0 = {1{$random}};
    seqLevelDoneReg2 = {1{$random}};
    bankSeqReg_0 = {3{$random}};
    bankSeqReg_1 = {3{$random}};
    bankSeqReg_2 = {3{$random}};
    bankSeqReg_3 = {3{$random}};
    bankSeqReg_4 = {3{$random}};
    bankSeqReg_5 = {3{$random}};
    bankSeqReg_6 = {3{$random}};
    bankSeqReg_7 = {3{$random}};
    seqLevelDoneReg1 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1 = T267 ? isReadValid : 1'h0;
  assign isReadValid = T2;
  assign T2 = T266 ? 1'h0 : T3;
  assign T3 = T267 ? localStorage_io_isReadValid_7 : T4;
  assign T4 = T265 ? 1'h0 : T5;
  assign T5 = T264 ? localStorage_io_isReadValid_6 : T6;
  assign T6 = T263 ? 1'h0 : T7;
  assign T7 = T262 ? localStorage_io_isReadValid_5 : T8;
  assign T8 = T261 ? 1'h0 : T9;
  assign T9 = T260 ? localStorage_io_isReadValid_4 : T10;
  assign T10 = T259 ? 1'h0 : T11;
  assign T11 = T258 ? localStorage_io_isReadValid_3 : T12;
  assign T12 = T257 ? 1'h0 : T13;
  assign T13 = T256 ? localStorage_io_isReadValid_2 : T14;
  assign T14 = T255 ? 1'h0 : T15;
  assign T15 = T254 ? localStorage_io_isReadValid_1 : T16;
  assign T16 = T17 ? localStorage_io_isReadValid_0 : 1'h0;
  assign T17 = T247 & T18;
  assign T18 = T19 & fifo_40_io_enqRdy;
  assign T19 = bankSeq[7'h57:7'h57];
  assign bankSeq = T20;
  assign T20 = T266 ? 88'h0 : T21;
  assign T21 = T240 ? T239 : T22;
  assign T22 = T265 ? 88'h0 : T23;
  assign T23 = T232 ? T231 : T24;
  assign T24 = T263 ? 88'h0 : T25;
  assign T25 = T224 ? T223 : T26;
  assign T26 = T261 ? 88'h0 : T27;
  assign T27 = T216 ? T215 : T28;
  assign T28 = T259 ? 88'h0 : T29;
  assign T29 = T208 ? T207 : T30;
  assign T30 = T257 ? 88'h0 : T31;
  assign T31 = T200 ? T199 : T32;
  assign T32 = T255 ? 88'h0 : T33;
  assign T33 = T183 ? T182 : T34;
  assign T34 = T247 ? T35 : 88'h0;
  assign T35 = nextSeq[7'h57:1'h0];
  assign nextSeq = T36;
  assign T36 = T266 ? 89'h0 : T37;
  assign T37 = T180 ? nextSeqReg2 : T38;
  assign T38 = T169 ? nextSeqReg2 : T39;
  assign T39 = T265 ? 89'h0 : T40;
  assign T40 = T167 ? nextSeqReg2 : T41;
  assign T41 = T166 ? nextSeqReg2 : T42;
  assign T42 = T263 ? 89'h0 : T43;
  assign T43 = T164 ? nextSeqReg2 : T44;
  assign T44 = T163 ? nextSeqReg2 : T45;
  assign T45 = T261 ? 89'h0 : T46;
  assign T46 = T161 ? nextSeqReg2 : T47;
  assign T47 = T160 ? nextSeqReg2 : T48;
  assign T48 = T259 ? 89'h0 : T49;
  assign T49 = T158 ? nextSeqReg2 : T50;
  assign T50 = T157 ? nextSeqReg2 : T51;
  assign T51 = T257 ? 89'h0 : T52;
  assign T52 = T155 ? nextSeqReg2 : T53;
  assign T53 = T154 ? nextSeqReg2 : T54;
  assign T54 = T255 ? 89'h0 : T55;
  assign T55 = T152 ? nextSeqReg2 : T56;
  assign T56 = T151 ? nextSeqReg2 : T57;
  assign T57 = T149 ? nextSeqReg2 : T58;
  assign T58 = T59 ? nextSeqReg2 : 89'h0;
  assign T59 = T247 & nextSeqSelReg;
  assign T3098 = reset ? 1'h0 : T60;
  assign T60 = fabInSeqMemConfig_io_rst ? 1'h0 : T61;
  assign T61 = allDone ? T62 : nextSeqSelReg;
  assign T62 = ~ nextSeqSelReg;
  assign allDone = T63;
  assign T63 = T74 & bankReadDone_7;
  assign bankReadDone_7 = T64;
  assign T64 = T266 ? 1'h0 : T65;
  assign T65 = T70 ? 1'h1 : T66;
  assign T66 = T68 ? 1'h0 : T67;
  assign T67 = T267 & isReadValid;
  assign T68 = T267 & T69;
  assign T69 = isReadValid ^ 1'h1;
  assign T70 = T240 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T73 & fifo_47_io_enqRdy;
  assign T73 = bankSeq[7'h57:7'h57];
  assign T74 = T85 & bankReadDone_6;
  assign bankReadDone_6 = T75;
  assign T75 = T265 ? 1'h0 : T76;
  assign T76 = T81 ? 1'h1 : T77;
  assign T77 = T79 ? 1'h0 : T78;
  assign T78 = T264 & isReadValid;
  assign T79 = T264 & T80;
  assign T80 = isReadValid ^ 1'h1;
  assign T81 = T232 & T82;
  assign T82 = T83 ^ 1'h1;
  assign T83 = T84 & fifo_46_io_enqRdy;
  assign T84 = bankSeq[7'h57:7'h57];
  assign T85 = T96 & bankReadDone_5;
  assign bankReadDone_5 = T86;
  assign T86 = T263 ? 1'h0 : T87;
  assign T87 = T92 ? 1'h1 : T88;
  assign T88 = T90 ? 1'h0 : T89;
  assign T89 = T262 & isReadValid;
  assign T90 = T262 & T91;
  assign T91 = isReadValid ^ 1'h1;
  assign T92 = T224 & T93;
  assign T93 = T94 ^ 1'h1;
  assign T94 = T95 & fifo_45_io_enqRdy;
  assign T95 = bankSeq[7'h57:7'h57];
  assign T96 = T107 & bankReadDone_4;
  assign bankReadDone_4 = T97;
  assign T97 = T261 ? 1'h0 : T98;
  assign T98 = T103 ? 1'h1 : T99;
  assign T99 = T101 ? 1'h0 : T100;
  assign T100 = T260 & isReadValid;
  assign T101 = T260 & T102;
  assign T102 = isReadValid ^ 1'h1;
  assign T103 = T216 & T104;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T106 & fifo_44_io_enqRdy;
  assign T106 = bankSeq[7'h57:7'h57];
  assign T107 = T118 & bankReadDone_3;
  assign bankReadDone_3 = T108;
  assign T108 = T259 ? 1'h0 : T109;
  assign T109 = T114 ? 1'h1 : T110;
  assign T110 = T112 ? 1'h0 : T111;
  assign T111 = T258 & isReadValid;
  assign T112 = T258 & T113;
  assign T113 = isReadValid ^ 1'h1;
  assign T114 = T208 & T115;
  assign T115 = T116 ^ 1'h1;
  assign T116 = T117 & fifo_43_io_enqRdy;
  assign T117 = bankSeq[7'h57:7'h57];
  assign T118 = T129 & bankReadDone_2;
  assign bankReadDone_2 = T119;
  assign T119 = T257 ? 1'h0 : T120;
  assign T120 = T125 ? 1'h1 : T121;
  assign T121 = T123 ? 1'h0 : T122;
  assign T122 = T256 & isReadValid;
  assign T123 = T256 & T124;
  assign T124 = isReadValid ^ 1'h1;
  assign T125 = T200 & T126;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T128 & fifo_42_io_enqRdy;
  assign T128 = bankSeq[7'h57:7'h57];
  assign T129 = bankReadDone_0 & bankReadDone_1;
  assign bankReadDone_1 = T130;
  assign T130 = T255 ? 1'h0 : T131;
  assign T131 = T136 ? 1'h1 : T132;
  assign T132 = T134 ? 1'h0 : T133;
  assign T133 = T254 & isReadValid;
  assign T134 = T254 & T135;
  assign T135 = isReadValid ^ 1'h1;
  assign T136 = T183 & T137;
  assign T137 = T138 ^ 1'h1;
  assign T138 = T139 & fifo_41_io_enqRdy;
  assign T139 = bankSeq[7'h57:7'h57];
  assign bankReadDone_0 = T140;
  assign T140 = T148 ? 1'h0 : T141;
  assign T141 = T146 ? 1'h1 : T142;
  assign T142 = T144 ? 1'h0 : T143;
  assign T143 = T17 & isReadValid;
  assign T144 = T17 & T145;
  assign T145 = isReadValid ^ 1'h1;
  assign T146 = T247 & T147;
  assign T147 = T18 ^ 1'h1;
  assign T148 = T247 ^ 1'h1;
  assign T149 = T247 & T150;
  assign T150 = nextSeqSelReg ^ 1'h1;
  assign T151 = T183 & nextSeqSelReg;
  assign T152 = T183 & T153;
  assign T153 = nextSeqSelReg ^ 1'h1;
  assign T154 = T200 & nextSeqSelReg;
  assign T155 = T200 & T156;
  assign T156 = nextSeqSelReg ^ 1'h1;
  assign T157 = T208 & nextSeqSelReg;
  assign T158 = T208 & T159;
  assign T159 = nextSeqSelReg ^ 1'h1;
  assign T160 = T216 & nextSeqSelReg;
  assign T161 = T216 & T162;
  assign T162 = nextSeqSelReg ^ 1'h1;
  assign T163 = T224 & nextSeqSelReg;
  assign T164 = T224 & T165;
  assign T165 = nextSeqSelReg ^ 1'h1;
  assign T166 = T232 & nextSeqSelReg;
  assign T167 = T232 & T168;
  assign T168 = nextSeqSelReg ^ 1'h1;
  assign T169 = T240 & nextSeqSelReg;
  assign T3099 = reset ? 89'h0 : T170;
  assign T170 = T174 ? nextSeqWire : nextSeqReg2;
  assign nextSeqWire = T171;
  assign T171 = T173 ? 89'h0 : T172;
  assign T172 = io_seqMemAddrValid ? fabInSeqMem_io_outData : 89'h0;
  assign T173 = io_seqMemAddrValid ^ 1'h1;
  assign T174 = T179 & firstSeqSelReg;
  assign T3100 = reset ? 1'h0 : T175;
  assign T175 = fabInSeqMemConfig_io_rst ? 1'h0 : T176;
  assign T176 = T177 ? 1'h1 : firstSeqSelReg;
  assign T177 = nextSeqSelReg | T178;
  assign T178 = ~ firstSeqSelReg;
  assign T179 = ~ nextSeqSelReg;
  assign T180 = T240 & T181;
  assign T181 = nextSeqSelReg ^ 1'h1;
  assign T182 = nextSeq[7'h57:1'h0];
  assign T183 = T189 & bankReadDoneReg_1;
  assign T3101 = reset ? 1'h0 : T184;
  assign T184 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_1;
  assign readDone_1 = T185;
  assign T185 = allDone ? 1'h0 : T186;
  assign T186 = T188 ? bankReadDoneReg_1 : T187;
  assign T187 = bankReadDone_1 ? 1'h1 : bankReadDoneReg_1;
  assign T188 = bankReadDone_1 ^ 1'h1;
  assign T189 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T3102 = reset ? 1'h0 : T190;
  assign T190 = fabInSeqMemConfig_io_rst ? 1'h0 : T191;
  assign T191 = T195 ? 1'h0 : T192;
  assign T192 = T194 ? 1'h0 : T193;
  assign T193 = T174 ? 1'h1 : nextSeqRegValid2;
  assign T194 = allDone & nextSeqSelReg;
  assign T195 = allDone & T196;
  assign T196 = nextSeqSelReg ^ 1'h1;
  assign T3103 = reset ? 1'h0 : T197;
  assign T197 = fabInSeqMemConfig_io_rst ? 1'h0 : T198;
  assign T198 = T177 ? 1'h1 : nextSeqRegValid1;
  assign T199 = nextSeq[7'h57:1'h0];
  assign T200 = T206 & bankReadDoneReg_2;
  assign T3104 = reset ? 1'h0 : T201;
  assign T201 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_2;
  assign readDone_2 = T202;
  assign T202 = allDone ? 1'h0 : T203;
  assign T203 = T205 ? bankReadDoneReg_2 : T204;
  assign T204 = bankReadDone_2 ? 1'h1 : bankReadDoneReg_2;
  assign T205 = bankReadDone_2 ^ 1'h1;
  assign T206 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T207 = nextSeq[7'h57:1'h0];
  assign T208 = T214 & bankReadDoneReg_3;
  assign T3105 = reset ? 1'h0 : T209;
  assign T209 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_3;
  assign readDone_3 = T210;
  assign T210 = allDone ? 1'h0 : T211;
  assign T211 = T213 ? bankReadDoneReg_3 : T212;
  assign T212 = bankReadDone_3 ? 1'h1 : bankReadDoneReg_3;
  assign T213 = bankReadDone_3 ^ 1'h1;
  assign T214 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T215 = nextSeq[7'h57:1'h0];
  assign T216 = T222 & bankReadDoneReg_4;
  assign T3106 = reset ? 1'h0 : T217;
  assign T217 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_4;
  assign readDone_4 = T218;
  assign T218 = allDone ? 1'h0 : T219;
  assign T219 = T221 ? bankReadDoneReg_4 : T220;
  assign T220 = bankReadDone_4 ? 1'h1 : bankReadDoneReg_4;
  assign T221 = bankReadDone_4 ^ 1'h1;
  assign T222 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T223 = nextSeq[7'h57:1'h0];
  assign T224 = T230 & bankReadDoneReg_5;
  assign T3107 = reset ? 1'h0 : T225;
  assign T225 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_5;
  assign readDone_5 = T226;
  assign T226 = allDone ? 1'h0 : T227;
  assign T227 = T229 ? bankReadDoneReg_5 : T228;
  assign T228 = bankReadDone_5 ? 1'h1 : bankReadDoneReg_5;
  assign T229 = bankReadDone_5 ^ 1'h1;
  assign T230 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T231 = nextSeq[7'h57:1'h0];
  assign T232 = T238 & bankReadDoneReg_6;
  assign T3108 = reset ? 1'h0 : T233;
  assign T233 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_6;
  assign readDone_6 = T234;
  assign T234 = allDone ? 1'h0 : T235;
  assign T235 = T237 ? bankReadDoneReg_6 : T236;
  assign T236 = bankReadDone_6 ? 1'h1 : bankReadDoneReg_6;
  assign T237 = bankReadDone_6 ^ 1'h1;
  assign T238 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T239 = nextSeq[7'h57:1'h0];
  assign T240 = T246 & bankReadDoneReg_7;
  assign T3109 = reset ? 1'h0 : T241;
  assign T241 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_7;
  assign readDone_7 = T242;
  assign T242 = allDone ? 1'h0 : T243;
  assign T243 = T245 ? bankReadDoneReg_7 : T244;
  assign T244 = bankReadDone_7 ? 1'h1 : bankReadDoneReg_7;
  assign T245 = bankReadDone_7 ^ 1'h1;
  assign T246 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T247 = T253 & bankReadDoneReg_0;
  assign T3110 = reset ? 1'h0 : T248;
  assign T248 = fabInSeqMemConfig_io_rst ? 1'h0 : readDone_0;
  assign readDone_0 = T249;
  assign T249 = allDone ? 1'h0 : T250;
  assign T250 = T252 ? bankReadDoneReg_0 : T251;
  assign T251 = bankReadDone_0 ? 1'h1 : bankReadDoneReg_0;
  assign T252 = bankReadDone_0 ^ 1'h1;
  assign T253 = nextSeqRegValid1 | nextSeqRegValid2;
  assign T254 = T183 & T138;
  assign T255 = T183 ^ 1'h1;
  assign T256 = T200 & T127;
  assign T257 = T200 ^ 1'h1;
  assign T258 = T208 & T116;
  assign T259 = T208 ^ 1'h1;
  assign T260 = T216 & T105;
  assign T261 = T216 ^ 1'h1;
  assign T262 = T224 & T94;
  assign T263 = T224 ^ 1'h1;
  assign T264 = T232 & T83;
  assign T265 = T232 ^ 1'h1;
  assign T266 = T240 ^ 1'h1;
  assign T267 = T240 & T72;
  assign T268 = T269 ? 1'h1 : 1'h0;
  assign T269 = T1568 | collectRdy;
  assign collectRdy = T270;
  assign T270 = T1567 ? 1'h0 : T271;
  assign T271 = T1565 ? 1'h0 : T272;
  assign T272 = seqLevelDoneReg2 & rdy;
  assign rdy = T273;
  assign T273 = seqLevelDoneReg2 ? T274 : 1'h0;
  assign T274 = rdyInit & T275;
  assign T275 = T277 & enqRdyCollect_19;
  assign enqRdyCollect_19 = T276;
  assign T276 = seqLevelDoneReg2 ? fifo_39_io_enqRdy : fifo_39_io_enqRdy;
  assign T277 = T279 & enqRdyCollect_18;
  assign enqRdyCollect_18 = T278;
  assign T278 = seqLevelDoneReg2 ? fifo_38_io_enqRdy : fifo_38_io_enqRdy;
  assign T279 = T281 & enqRdyCollect_17;
  assign enqRdyCollect_17 = T280;
  assign T280 = seqLevelDoneReg2 ? fifo_37_io_enqRdy : fifo_37_io_enqRdy;
  assign T281 = T283 & enqRdyCollect_16;
  assign enqRdyCollect_16 = T282;
  assign T282 = seqLevelDoneReg2 ? fifo_36_io_enqRdy : fifo_36_io_enqRdy;
  assign T283 = T285 & enqRdyCollect_15;
  assign enqRdyCollect_15 = T284;
  assign T284 = seqLevelDoneReg2 ? fifo_35_io_enqRdy : fifo_35_io_enqRdy;
  assign T285 = T287 & enqRdyCollect_14;
  assign enqRdyCollect_14 = T286;
  assign T286 = seqLevelDoneReg2 ? fifo_34_io_enqRdy : fifo_34_io_enqRdy;
  assign T287 = T289 & enqRdyCollect_13;
  assign enqRdyCollect_13 = T288;
  assign T288 = seqLevelDoneReg2 ? fifo_33_io_enqRdy : fifo_33_io_enqRdy;
  assign T289 = T291 & enqRdyCollect_12;
  assign enqRdyCollect_12 = T290;
  assign T290 = seqLevelDoneReg2 ? fifo_32_io_enqRdy : fifo_32_io_enqRdy;
  assign T291 = T293 & enqRdyCollect_11;
  assign enqRdyCollect_11 = T292;
  assign T292 = seqLevelDoneReg2 ? fifo_31_io_enqRdy : fifo_31_io_enqRdy;
  assign T293 = T295 & enqRdyCollect_10;
  assign enqRdyCollect_10 = T294;
  assign T294 = seqLevelDoneReg2 ? fifo_30_io_enqRdy : fifo_30_io_enqRdy;
  assign T295 = T297 & enqRdyCollect_9;
  assign enqRdyCollect_9 = T296;
  assign T296 = seqLevelDoneReg2 ? fifo_29_io_enqRdy : fifo_29_io_enqRdy;
  assign T297 = T299 & enqRdyCollect_8;
  assign enqRdyCollect_8 = T298;
  assign T298 = seqLevelDoneReg2 ? fifo_28_io_enqRdy : fifo_28_io_enqRdy;
  assign T299 = T301 & enqRdyCollect_7;
  assign enqRdyCollect_7 = T300;
  assign T300 = seqLevelDoneReg2 ? fifo_27_io_enqRdy : fifo_27_io_enqRdy;
  assign T301 = T303 & enqRdyCollect_6;
  assign enqRdyCollect_6 = T302;
  assign T302 = seqLevelDoneReg2 ? fifo_26_io_enqRdy : fifo_26_io_enqRdy;
  assign T303 = T305 & enqRdyCollect_5;
  assign enqRdyCollect_5 = T304;
  assign T304 = seqLevelDoneReg2 ? fifo_25_io_enqRdy : fifo_25_io_enqRdy;
  assign T305 = T307 & enqRdyCollect_4;
  assign enqRdyCollect_4 = T306;
  assign T306 = seqLevelDoneReg2 ? fifo_24_io_enqRdy : fifo_24_io_enqRdy;
  assign T307 = T309 & enqRdyCollect_3;
  assign enqRdyCollect_3 = T308;
  assign T308 = seqLevelDoneReg2 ? fifo_23_io_enqRdy : fifo_23_io_enqRdy;
  assign T309 = T311 & enqRdyCollect_2;
  assign enqRdyCollect_2 = T310;
  assign T310 = seqLevelDoneReg2 ? fifo_22_io_enqRdy : fifo_22_io_enqRdy;
  assign T311 = enqRdyCollect_0 & enqRdyCollect_1;
  assign enqRdyCollect_1 = T312;
  assign T312 = seqLevelDoneReg2 ? fifo_21_io_enqRdy : fifo_21_io_enqRdy;
  assign enqRdyCollect_0 = T313;
  assign T313 = seqLevelDoneReg2 ? fifo_20_io_enqRdy : fifo_20_io_enqRdy;
  assign rdyInit = T314;
  assign T314 = seqLevelDoneReg2 ? 1'h1 : 1'h0;
  assign T3111 = reset ? 1'h0 : T315;
  assign T315 = fabInSeqMemConfig_io_rst ? 1'h0 : T316;
  assign T316 = T1509 ? seqLevelDoneReg1 : T317;
  assign T317 = T1453 ? seqLevelDoneReg1 : T318;
  assign T318 = T1397 ? seqLevelDoneReg1 : T319;
  assign T319 = T1341 ? seqLevelDoneReg1 : T320;
  assign T320 = T1285 ? seqLevelDoneReg1 : T321;
  assign T321 = T1229 ? seqLevelDoneReg1 : T322;
  assign T322 = T1173 ? seqLevelDoneReg1 : T323;
  assign T323 = T1117 ? seqLevelDoneReg1 : T324;
  assign T324 = T1061 ? seqLevelDoneReg1 : T325;
  assign T325 = T1005 ? seqLevelDoneReg1 : T326;
  assign T326 = T949 ? seqLevelDoneReg1 : T327;
  assign T327 = T893 ? seqLevelDoneReg1 : T328;
  assign T328 = T837 ? seqLevelDoneReg1 : T329;
  assign T329 = T781 ? seqLevelDoneReg1 : T330;
  assign T330 = T725 ? seqLevelDoneReg1 : T331;
  assign T331 = T669 ? seqLevelDoneReg1 : T332;
  assign T332 = T613 ? seqLevelDoneReg1 : T333;
  assign T333 = T557 ? seqLevelDoneReg1 : T334;
  assign T334 = T501 ? seqLevelDoneReg1 : T335;
  assign T335 = T361 ? seqLevelDoneReg1 : seqLevelDoneReg2;
  assign T361 = T362;
  assign T362 = T438 & T363;
  assign T363 = bankToPortValid_7_0;
  assign bankToPortValid_7_0 = T364;
  assign T364 = T437 ? 1'h0 : T365;
  assign T365 = T366 ? fifo_47_io_deqValid : 1'h0;
  assign T366 = T269 & T367;
  assign T367 = T368[1'h0:1'h0];
  assign T368 = 1'h1 << T369;
  assign T369 = T3112;
  assign T3112 = {2'h0, portId};
  assign portId = T370;
  assign T370 = T436 ? T435 : T371;
  assign T371 = T269 ? T434 : T372;
  assign T372 = T433 ? T432 : T373;
  assign T373 = T430 ? T429 : T374;
  assign T374 = T428 ? T427 : T375;
  assign T375 = T425 ? T424 : T376;
  assign T376 = T423 ? T422 : T377;
  assign T377 = T420 ? T419 : T378;
  assign T378 = T418 ? T417 : T379;
  assign T379 = T415 ? T414 : T380;
  assign T380 = T413 ? T412 : T381;
  assign T381 = T410 ? T409 : T382;
  assign T382 = T408 ? T407 : T383;
  assign T383 = T405 ? T404 : T384;
  assign T384 = T402 ? T401 : T385;
  assign T385 = bankSeq2[2'h2:1'h0];
  assign bankSeq2 = T386;
  assign T386 = T436 ? bankSeqReg_7 : T387;
  assign T387 = T269 ? bankSeqReg_7 : T388;
  assign T388 = T433 ? bankSeqReg_6 : T389;
  assign T389 = T430 ? bankSeqReg_6 : T390;
  assign T390 = T428 ? bankSeqReg_5 : T391;
  assign T391 = T425 ? bankSeqReg_5 : T392;
  assign T392 = T423 ? bankSeqReg_4 : T393;
  assign T393 = T420 ? bankSeqReg_4 : T394;
  assign T394 = T418 ? bankSeqReg_3 : T395;
  assign T395 = T415 ? bankSeqReg_3 : T396;
  assign T396 = T413 ? bankSeqReg_2 : T397;
  assign T397 = T410 ? bankSeqReg_2 : T398;
  assign T398 = T408 ? bankSeqReg_1 : T399;
  assign T399 = T405 ? bankSeqReg_1 : T400;
  assign T400 = T402 ? bankSeqReg_0 : bankSeqReg_0;
  assign T3113 = reset ? 88'h0 : bankSeqReg_0;
  assign T3114 = reset ? 88'h0 : bankSeqReg_1;
  assign T3115 = reset ? 88'h0 : bankSeqReg_2;
  assign T3116 = reset ? 88'h0 : bankSeqReg_3;
  assign T3117 = reset ? 88'h0 : bankSeqReg_4;
  assign T3118 = reset ? 88'h0 : bankSeqReg_5;
  assign T3119 = reset ? 88'h0 : bankSeqReg_6;
  assign T3120 = reset ? 88'h0 : bankSeqReg_7;
  assign T401 = bankSeq2[2'h2:1'h0];
  assign T402 = T403 | collectRdy;
  assign T403 = ~ seqLevelDoneReg2;
  assign T404 = bankSeq2[2'h2:1'h0];
  assign T405 = T406 | collectRdy;
  assign T406 = ~ seqLevelDoneReg2;
  assign T407 = bankSeq2[2'h2:1'h0];
  assign T408 = T405 ^ 1'h1;
  assign T409 = bankSeq2[2'h2:1'h0];
  assign T410 = T411 | collectRdy;
  assign T411 = ~ seqLevelDoneReg2;
  assign T412 = bankSeq2[2'h2:1'h0];
  assign T413 = T410 ^ 1'h1;
  assign T414 = bankSeq2[2'h2:1'h0];
  assign T415 = T416 | collectRdy;
  assign T416 = ~ seqLevelDoneReg2;
  assign T417 = bankSeq2[2'h2:1'h0];
  assign T418 = T415 ^ 1'h1;
  assign T419 = bankSeq2[2'h2:1'h0];
  assign T420 = T421 | collectRdy;
  assign T421 = ~ seqLevelDoneReg2;
  assign T422 = bankSeq2[2'h2:1'h0];
  assign T423 = T420 ^ 1'h1;
  assign T424 = bankSeq2[2'h2:1'h0];
  assign T425 = T426 | collectRdy;
  assign T426 = ~ seqLevelDoneReg2;
  assign T427 = bankSeq2[2'h2:1'h0];
  assign T428 = T425 ^ 1'h1;
  assign T429 = bankSeq2[2'h2:1'h0];
  assign T430 = T431 | collectRdy;
  assign T431 = ~ seqLevelDoneReg2;
  assign T432 = bankSeq2[2'h2:1'h0];
  assign T433 = T430 ^ 1'h1;
  assign T434 = bankSeq2[2'h2:1'h0];
  assign T435 = bankSeq2[2'h2:1'h0];
  assign T436 = T269 ^ 1'h1;
  assign T437 = T436 & T367;
  assign T438 = T447 & T439;
  assign T439 = bankToPortValid_6_0;
  assign bankToPortValid_6_0 = T440;
  assign T440 = T446 ? 1'h0 : T441;
  assign T441 = T442 ? fifo_46_io_deqValid : 1'h0;
  assign T442 = T430 & T443;
  assign T443 = T444[1'h0:1'h0];
  assign T444 = 1'h1 << T445;
  assign T445 = T3121;
  assign T3121 = {2'h0, portId};
  assign T446 = T433 & T443;
  assign T447 = T456 & T448;
  assign T448 = bankToPortValid_5_0;
  assign bankToPortValid_5_0 = T449;
  assign T449 = T455 ? 1'h0 : T450;
  assign T450 = T451 ? fifo_45_io_deqValid : 1'h0;
  assign T451 = T425 & T452;
  assign T452 = T453[1'h0:1'h0];
  assign T453 = 1'h1 << T454;
  assign T454 = T3122;
  assign T3122 = {2'h0, portId};
  assign T455 = T428 & T452;
  assign T456 = T465 & T457;
  assign T457 = bankToPortValid_4_0;
  assign bankToPortValid_4_0 = T458;
  assign T458 = T464 ? 1'h0 : T459;
  assign T459 = T460 ? fifo_44_io_deqValid : 1'h0;
  assign T460 = T420 & T461;
  assign T461 = T462[1'h0:1'h0];
  assign T462 = 1'h1 << T463;
  assign T463 = T3123;
  assign T3123 = {2'h0, portId};
  assign T464 = T423 & T461;
  assign T465 = T474 & T466;
  assign T466 = bankToPortValid_3_0;
  assign bankToPortValid_3_0 = T467;
  assign T467 = T473 ? 1'h0 : T468;
  assign T468 = T469 ? fifo_43_io_deqValid : 1'h0;
  assign T469 = T415 & T470;
  assign T470 = T471[1'h0:1'h0];
  assign T471 = 1'h1 << T472;
  assign T472 = T3124;
  assign T3124 = {2'h0, portId};
  assign T473 = T418 & T470;
  assign T474 = T483 & T475;
  assign T475 = bankToPortValid_2_0;
  assign bankToPortValid_2_0 = T476;
  assign T476 = T482 ? 1'h0 : T477;
  assign T477 = T478 ? fifo_42_io_deqValid : 1'h0;
  assign T478 = T410 & T479;
  assign T479 = T480[1'h0:1'h0];
  assign T480 = 1'h1 << T481;
  assign T481 = T3125;
  assign T3125 = {2'h0, portId};
  assign T482 = T413 & T479;
  assign T483 = T492 & T484;
  assign T484 = bankToPortValid_1_0;
  assign bankToPortValid_1_0 = T485;
  assign T485 = T491 ? 1'h0 : T486;
  assign T486 = T487 ? fifo_41_io_deqValid : 1'h0;
  assign T487 = T405 & T488;
  assign T488 = T489[1'h0:1'h0];
  assign T489 = 1'h1 << T490;
  assign T490 = T3126;
  assign T3126 = {2'h0, portId};
  assign T491 = T408 & T488;
  assign T492 = bankToPortValid_0_0;
  assign bankToPortValid_0_0 = T493;
  assign T493 = T499 ? 1'h0 : T494;
  assign T494 = T495 ? fifo_40_io_deqValid : 1'h0;
  assign T495 = T402 & T496;
  assign T496 = T497[1'h0:1'h0];
  assign T497 = 1'h1 << T498;
  assign T498 = T3127;
  assign T3127 = {2'h0, portId};
  assign T499 = T500 & T496;
  assign T500 = T402 ^ 1'h1;
  assign T501 = T502;
  assign T502 = T509 & T503;
  assign T503 = bankToPortValid_7_1;
  assign bankToPortValid_7_1 = T504;
  assign T504 = T508 ? 1'h0 : T505;
  assign T505 = T506 ? fifo_47_io_deqValid : 1'h0;
  assign T506 = T269 & T507;
  assign T507 = T368[1'h1:1'h1];
  assign T508 = T436 & T507;
  assign T509 = T516 & T510;
  assign T510 = bankToPortValid_6_1;
  assign bankToPortValid_6_1 = T511;
  assign T511 = T515 ? 1'h0 : T512;
  assign T512 = T513 ? fifo_46_io_deqValid : 1'h0;
  assign T513 = T430 & T514;
  assign T514 = T444[1'h1:1'h1];
  assign T515 = T433 & T514;
  assign T516 = T523 & T517;
  assign T517 = bankToPortValid_5_1;
  assign bankToPortValid_5_1 = T518;
  assign T518 = T522 ? 1'h0 : T519;
  assign T519 = T520 ? fifo_45_io_deqValid : 1'h0;
  assign T520 = T425 & T521;
  assign T521 = T453[1'h1:1'h1];
  assign T522 = T428 & T521;
  assign T523 = T530 & T524;
  assign T524 = bankToPortValid_4_1;
  assign bankToPortValid_4_1 = T525;
  assign T525 = T529 ? 1'h0 : T526;
  assign T526 = T527 ? fifo_44_io_deqValid : 1'h0;
  assign T527 = T420 & T528;
  assign T528 = T462[1'h1:1'h1];
  assign T529 = T423 & T528;
  assign T530 = T537 & T531;
  assign T531 = bankToPortValid_3_1;
  assign bankToPortValid_3_1 = T532;
  assign T532 = T536 ? 1'h0 : T533;
  assign T533 = T534 ? fifo_43_io_deqValid : 1'h0;
  assign T534 = T415 & T535;
  assign T535 = T471[1'h1:1'h1];
  assign T536 = T418 & T535;
  assign T537 = T544 & T538;
  assign T538 = bankToPortValid_2_1;
  assign bankToPortValid_2_1 = T539;
  assign T539 = T543 ? 1'h0 : T540;
  assign T540 = T541 ? fifo_42_io_deqValid : 1'h0;
  assign T541 = T410 & T542;
  assign T542 = T480[1'h1:1'h1];
  assign T543 = T413 & T542;
  assign T544 = T551 & T545;
  assign T545 = bankToPortValid_1_1;
  assign bankToPortValid_1_1 = T546;
  assign T546 = T550 ? 1'h0 : T547;
  assign T547 = T548 ? fifo_41_io_deqValid : 1'h0;
  assign T548 = T405 & T549;
  assign T549 = T489[1'h1:1'h1];
  assign T550 = T408 & T549;
  assign T551 = bankToPortValid_0_1;
  assign bankToPortValid_0_1 = T552;
  assign T552 = T556 ? 1'h0 : T553;
  assign T553 = T554 ? fifo_40_io_deqValid : 1'h0;
  assign T554 = T402 & T555;
  assign T555 = T497[1'h1:1'h1];
  assign T556 = T500 & T555;
  assign T557 = T558;
  assign T558 = T565 & T559;
  assign T559 = bankToPortValid_7_2;
  assign bankToPortValid_7_2 = T560;
  assign T560 = T564 ? 1'h0 : T561;
  assign T561 = T562 ? fifo_47_io_deqValid : 1'h0;
  assign T562 = T269 & T563;
  assign T563 = T368[2'h2:2'h2];
  assign T564 = T436 & T563;
  assign T565 = T572 & T566;
  assign T566 = bankToPortValid_6_2;
  assign bankToPortValid_6_2 = T567;
  assign T567 = T571 ? 1'h0 : T568;
  assign T568 = T569 ? fifo_46_io_deqValid : 1'h0;
  assign T569 = T430 & T570;
  assign T570 = T444[2'h2:2'h2];
  assign T571 = T433 & T570;
  assign T572 = T579 & T573;
  assign T573 = bankToPortValid_5_2;
  assign bankToPortValid_5_2 = T574;
  assign T574 = T578 ? 1'h0 : T575;
  assign T575 = T576 ? fifo_45_io_deqValid : 1'h0;
  assign T576 = T425 & T577;
  assign T577 = T453[2'h2:2'h2];
  assign T578 = T428 & T577;
  assign T579 = T586 & T580;
  assign T580 = bankToPortValid_4_2;
  assign bankToPortValid_4_2 = T581;
  assign T581 = T585 ? 1'h0 : T582;
  assign T582 = T583 ? fifo_44_io_deqValid : 1'h0;
  assign T583 = T420 & T584;
  assign T584 = T462[2'h2:2'h2];
  assign T585 = T423 & T584;
  assign T586 = T593 & T587;
  assign T587 = bankToPortValid_3_2;
  assign bankToPortValid_3_2 = T588;
  assign T588 = T592 ? 1'h0 : T589;
  assign T589 = T590 ? fifo_43_io_deqValid : 1'h0;
  assign T590 = T415 & T591;
  assign T591 = T471[2'h2:2'h2];
  assign T592 = T418 & T591;
  assign T593 = T600 & T594;
  assign T594 = bankToPortValid_2_2;
  assign bankToPortValid_2_2 = T595;
  assign T595 = T599 ? 1'h0 : T596;
  assign T596 = T597 ? fifo_42_io_deqValid : 1'h0;
  assign T597 = T410 & T598;
  assign T598 = T480[2'h2:2'h2];
  assign T599 = T413 & T598;
  assign T600 = T607 & T601;
  assign T601 = bankToPortValid_1_2;
  assign bankToPortValid_1_2 = T602;
  assign T602 = T606 ? 1'h0 : T603;
  assign T603 = T604 ? fifo_41_io_deqValid : 1'h0;
  assign T604 = T405 & T605;
  assign T605 = T489[2'h2:2'h2];
  assign T606 = T408 & T605;
  assign T607 = bankToPortValid_0_2;
  assign bankToPortValid_0_2 = T608;
  assign T608 = T612 ? 1'h0 : T609;
  assign T609 = T610 ? fifo_40_io_deqValid : 1'h0;
  assign T610 = T402 & T611;
  assign T611 = T497[2'h2:2'h2];
  assign T612 = T500 & T611;
  assign T613 = T614;
  assign T614 = T621 & T615;
  assign T615 = bankToPortValid_7_3;
  assign bankToPortValid_7_3 = T616;
  assign T616 = T620 ? 1'h0 : T617;
  assign T617 = T618 ? fifo_47_io_deqValid : 1'h0;
  assign T618 = T269 & T619;
  assign T619 = T368[2'h3:2'h3];
  assign T620 = T436 & T619;
  assign T621 = T628 & T622;
  assign T622 = bankToPortValid_6_3;
  assign bankToPortValid_6_3 = T623;
  assign T623 = T627 ? 1'h0 : T624;
  assign T624 = T625 ? fifo_46_io_deqValid : 1'h0;
  assign T625 = T430 & T626;
  assign T626 = T444[2'h3:2'h3];
  assign T627 = T433 & T626;
  assign T628 = T635 & T629;
  assign T629 = bankToPortValid_5_3;
  assign bankToPortValid_5_3 = T630;
  assign T630 = T634 ? 1'h0 : T631;
  assign T631 = T632 ? fifo_45_io_deqValid : 1'h0;
  assign T632 = T425 & T633;
  assign T633 = T453[2'h3:2'h3];
  assign T634 = T428 & T633;
  assign T635 = T642 & T636;
  assign T636 = bankToPortValid_4_3;
  assign bankToPortValid_4_3 = T637;
  assign T637 = T641 ? 1'h0 : T638;
  assign T638 = T639 ? fifo_44_io_deqValid : 1'h0;
  assign T639 = T420 & T640;
  assign T640 = T462[2'h3:2'h3];
  assign T641 = T423 & T640;
  assign T642 = T649 & T643;
  assign T643 = bankToPortValid_3_3;
  assign bankToPortValid_3_3 = T644;
  assign T644 = T648 ? 1'h0 : T645;
  assign T645 = T646 ? fifo_43_io_deqValid : 1'h0;
  assign T646 = T415 & T647;
  assign T647 = T471[2'h3:2'h3];
  assign T648 = T418 & T647;
  assign T649 = T656 & T650;
  assign T650 = bankToPortValid_2_3;
  assign bankToPortValid_2_3 = T651;
  assign T651 = T655 ? 1'h0 : T652;
  assign T652 = T653 ? fifo_42_io_deqValid : 1'h0;
  assign T653 = T410 & T654;
  assign T654 = T480[2'h3:2'h3];
  assign T655 = T413 & T654;
  assign T656 = T663 & T657;
  assign T657 = bankToPortValid_1_3;
  assign bankToPortValid_1_3 = T658;
  assign T658 = T662 ? 1'h0 : T659;
  assign T659 = T660 ? fifo_41_io_deqValid : 1'h0;
  assign T660 = T405 & T661;
  assign T661 = T489[2'h3:2'h3];
  assign T662 = T408 & T661;
  assign T663 = bankToPortValid_0_3;
  assign bankToPortValid_0_3 = T664;
  assign T664 = T668 ? 1'h0 : T665;
  assign T665 = T666 ? fifo_40_io_deqValid : 1'h0;
  assign T666 = T402 & T667;
  assign T667 = T497[2'h3:2'h3];
  assign T668 = T500 & T667;
  assign T669 = T670;
  assign T670 = T677 & T671;
  assign T671 = bankToPortValid_7_4;
  assign bankToPortValid_7_4 = T672;
  assign T672 = T676 ? 1'h0 : T673;
  assign T673 = T674 ? fifo_47_io_deqValid : 1'h0;
  assign T674 = T269 & T675;
  assign T675 = T368[3'h4:3'h4];
  assign T676 = T436 & T675;
  assign T677 = T684 & T678;
  assign T678 = bankToPortValid_6_4;
  assign bankToPortValid_6_4 = T679;
  assign T679 = T683 ? 1'h0 : T680;
  assign T680 = T681 ? fifo_46_io_deqValid : 1'h0;
  assign T681 = T430 & T682;
  assign T682 = T444[3'h4:3'h4];
  assign T683 = T433 & T682;
  assign T684 = T691 & T685;
  assign T685 = bankToPortValid_5_4;
  assign bankToPortValid_5_4 = T686;
  assign T686 = T690 ? 1'h0 : T687;
  assign T687 = T688 ? fifo_45_io_deqValid : 1'h0;
  assign T688 = T425 & T689;
  assign T689 = T453[3'h4:3'h4];
  assign T690 = T428 & T689;
  assign T691 = T698 & T692;
  assign T692 = bankToPortValid_4_4;
  assign bankToPortValid_4_4 = T693;
  assign T693 = T697 ? 1'h0 : T694;
  assign T694 = T695 ? fifo_44_io_deqValid : 1'h0;
  assign T695 = T420 & T696;
  assign T696 = T462[3'h4:3'h4];
  assign T697 = T423 & T696;
  assign T698 = T705 & T699;
  assign T699 = bankToPortValid_3_4;
  assign bankToPortValid_3_4 = T700;
  assign T700 = T704 ? 1'h0 : T701;
  assign T701 = T702 ? fifo_43_io_deqValid : 1'h0;
  assign T702 = T415 & T703;
  assign T703 = T471[3'h4:3'h4];
  assign T704 = T418 & T703;
  assign T705 = T712 & T706;
  assign T706 = bankToPortValid_2_4;
  assign bankToPortValid_2_4 = T707;
  assign T707 = T711 ? 1'h0 : T708;
  assign T708 = T709 ? fifo_42_io_deqValid : 1'h0;
  assign T709 = T410 & T710;
  assign T710 = T480[3'h4:3'h4];
  assign T711 = T413 & T710;
  assign T712 = T719 & T713;
  assign T713 = bankToPortValid_1_4;
  assign bankToPortValid_1_4 = T714;
  assign T714 = T718 ? 1'h0 : T715;
  assign T715 = T716 ? fifo_41_io_deqValid : 1'h0;
  assign T716 = T405 & T717;
  assign T717 = T489[3'h4:3'h4];
  assign T718 = T408 & T717;
  assign T719 = bankToPortValid_0_4;
  assign bankToPortValid_0_4 = T720;
  assign T720 = T724 ? 1'h0 : T721;
  assign T721 = T722 ? fifo_40_io_deqValid : 1'h0;
  assign T722 = T402 & T723;
  assign T723 = T497[3'h4:3'h4];
  assign T724 = T500 & T723;
  assign T725 = T726;
  assign T726 = T733 & T727;
  assign T727 = bankToPortValid_7_5;
  assign bankToPortValid_7_5 = T728;
  assign T728 = T732 ? 1'h0 : T729;
  assign T729 = T730 ? fifo_47_io_deqValid : 1'h0;
  assign T730 = T269 & T731;
  assign T731 = T368[3'h5:3'h5];
  assign T732 = T436 & T731;
  assign T733 = T740 & T734;
  assign T734 = bankToPortValid_6_5;
  assign bankToPortValid_6_5 = T735;
  assign T735 = T739 ? 1'h0 : T736;
  assign T736 = T737 ? fifo_46_io_deqValid : 1'h0;
  assign T737 = T430 & T738;
  assign T738 = T444[3'h5:3'h5];
  assign T739 = T433 & T738;
  assign T740 = T747 & T741;
  assign T741 = bankToPortValid_5_5;
  assign bankToPortValid_5_5 = T742;
  assign T742 = T746 ? 1'h0 : T743;
  assign T743 = T744 ? fifo_45_io_deqValid : 1'h0;
  assign T744 = T425 & T745;
  assign T745 = T453[3'h5:3'h5];
  assign T746 = T428 & T745;
  assign T747 = T754 & T748;
  assign T748 = bankToPortValid_4_5;
  assign bankToPortValid_4_5 = T749;
  assign T749 = T753 ? 1'h0 : T750;
  assign T750 = T751 ? fifo_44_io_deqValid : 1'h0;
  assign T751 = T420 & T752;
  assign T752 = T462[3'h5:3'h5];
  assign T753 = T423 & T752;
  assign T754 = T761 & T755;
  assign T755 = bankToPortValid_3_5;
  assign bankToPortValid_3_5 = T756;
  assign T756 = T760 ? 1'h0 : T757;
  assign T757 = T758 ? fifo_43_io_deqValid : 1'h0;
  assign T758 = T415 & T759;
  assign T759 = T471[3'h5:3'h5];
  assign T760 = T418 & T759;
  assign T761 = T768 & T762;
  assign T762 = bankToPortValid_2_5;
  assign bankToPortValid_2_5 = T763;
  assign T763 = T767 ? 1'h0 : T764;
  assign T764 = T765 ? fifo_42_io_deqValid : 1'h0;
  assign T765 = T410 & T766;
  assign T766 = T480[3'h5:3'h5];
  assign T767 = T413 & T766;
  assign T768 = T775 & T769;
  assign T769 = bankToPortValid_1_5;
  assign bankToPortValid_1_5 = T770;
  assign T770 = T774 ? 1'h0 : T771;
  assign T771 = T772 ? fifo_41_io_deqValid : 1'h0;
  assign T772 = T405 & T773;
  assign T773 = T489[3'h5:3'h5];
  assign T774 = T408 & T773;
  assign T775 = bankToPortValid_0_5;
  assign bankToPortValid_0_5 = T776;
  assign T776 = T780 ? 1'h0 : T777;
  assign T777 = T778 ? fifo_40_io_deqValid : 1'h0;
  assign T778 = T402 & T779;
  assign T779 = T497[3'h5:3'h5];
  assign T780 = T500 & T779;
  assign T781 = T782;
  assign T782 = T789 & T783;
  assign T783 = bankToPortValid_7_6;
  assign bankToPortValid_7_6 = T784;
  assign T784 = T788 ? 1'h0 : T785;
  assign T785 = T786 ? fifo_47_io_deqValid : 1'h0;
  assign T786 = T269 & T787;
  assign T787 = T368[3'h6:3'h6];
  assign T788 = T436 & T787;
  assign T789 = T796 & T790;
  assign T790 = bankToPortValid_6_6;
  assign bankToPortValid_6_6 = T791;
  assign T791 = T795 ? 1'h0 : T792;
  assign T792 = T793 ? fifo_46_io_deqValid : 1'h0;
  assign T793 = T430 & T794;
  assign T794 = T444[3'h6:3'h6];
  assign T795 = T433 & T794;
  assign T796 = T803 & T797;
  assign T797 = bankToPortValid_5_6;
  assign bankToPortValid_5_6 = T798;
  assign T798 = T802 ? 1'h0 : T799;
  assign T799 = T800 ? fifo_45_io_deqValid : 1'h0;
  assign T800 = T425 & T801;
  assign T801 = T453[3'h6:3'h6];
  assign T802 = T428 & T801;
  assign T803 = T810 & T804;
  assign T804 = bankToPortValid_4_6;
  assign bankToPortValid_4_6 = T805;
  assign T805 = T809 ? 1'h0 : T806;
  assign T806 = T807 ? fifo_44_io_deqValid : 1'h0;
  assign T807 = T420 & T808;
  assign T808 = T462[3'h6:3'h6];
  assign T809 = T423 & T808;
  assign T810 = T817 & T811;
  assign T811 = bankToPortValid_3_6;
  assign bankToPortValid_3_6 = T812;
  assign T812 = T816 ? 1'h0 : T813;
  assign T813 = T814 ? fifo_43_io_deqValid : 1'h0;
  assign T814 = T415 & T815;
  assign T815 = T471[3'h6:3'h6];
  assign T816 = T418 & T815;
  assign T817 = T824 & T818;
  assign T818 = bankToPortValid_2_6;
  assign bankToPortValid_2_6 = T819;
  assign T819 = T823 ? 1'h0 : T820;
  assign T820 = T821 ? fifo_42_io_deqValid : 1'h0;
  assign T821 = T410 & T822;
  assign T822 = T480[3'h6:3'h6];
  assign T823 = T413 & T822;
  assign T824 = T831 & T825;
  assign T825 = bankToPortValid_1_6;
  assign bankToPortValid_1_6 = T826;
  assign T826 = T830 ? 1'h0 : T827;
  assign T827 = T828 ? fifo_41_io_deqValid : 1'h0;
  assign T828 = T405 & T829;
  assign T829 = T489[3'h6:3'h6];
  assign T830 = T408 & T829;
  assign T831 = bankToPortValid_0_6;
  assign bankToPortValid_0_6 = T832;
  assign T832 = T836 ? 1'h0 : T833;
  assign T833 = T834 ? fifo_40_io_deqValid : 1'h0;
  assign T834 = T402 & T835;
  assign T835 = T497[3'h6:3'h6];
  assign T836 = T500 & T835;
  assign T837 = T838;
  assign T838 = T845 & T839;
  assign T839 = bankToPortValid_7_7;
  assign bankToPortValid_7_7 = T840;
  assign T840 = T844 ? 1'h0 : T841;
  assign T841 = T842 ? fifo_47_io_deqValid : 1'h0;
  assign T842 = T269 & T843;
  assign T843 = T368[3'h7:3'h7];
  assign T844 = T436 & T843;
  assign T845 = T852 & T846;
  assign T846 = bankToPortValid_6_7;
  assign bankToPortValid_6_7 = T847;
  assign T847 = T851 ? 1'h0 : T848;
  assign T848 = T849 ? fifo_46_io_deqValid : 1'h0;
  assign T849 = T430 & T850;
  assign T850 = T444[3'h7:3'h7];
  assign T851 = T433 & T850;
  assign T852 = T859 & T853;
  assign T853 = bankToPortValid_5_7;
  assign bankToPortValid_5_7 = T854;
  assign T854 = T858 ? 1'h0 : T855;
  assign T855 = T856 ? fifo_45_io_deqValid : 1'h0;
  assign T856 = T425 & T857;
  assign T857 = T453[3'h7:3'h7];
  assign T858 = T428 & T857;
  assign T859 = T866 & T860;
  assign T860 = bankToPortValid_4_7;
  assign bankToPortValid_4_7 = T861;
  assign T861 = T865 ? 1'h0 : T862;
  assign T862 = T863 ? fifo_44_io_deqValid : 1'h0;
  assign T863 = T420 & T864;
  assign T864 = T462[3'h7:3'h7];
  assign T865 = T423 & T864;
  assign T866 = T873 & T867;
  assign T867 = bankToPortValid_3_7;
  assign bankToPortValid_3_7 = T868;
  assign T868 = T872 ? 1'h0 : T869;
  assign T869 = T870 ? fifo_43_io_deqValid : 1'h0;
  assign T870 = T415 & T871;
  assign T871 = T471[3'h7:3'h7];
  assign T872 = T418 & T871;
  assign T873 = T880 & T874;
  assign T874 = bankToPortValid_2_7;
  assign bankToPortValid_2_7 = T875;
  assign T875 = T879 ? 1'h0 : T876;
  assign T876 = T877 ? fifo_42_io_deqValid : 1'h0;
  assign T877 = T410 & T878;
  assign T878 = T480[3'h7:3'h7];
  assign T879 = T413 & T878;
  assign T880 = T887 & T881;
  assign T881 = bankToPortValid_1_7;
  assign bankToPortValid_1_7 = T882;
  assign T882 = T886 ? 1'h0 : T883;
  assign T883 = T884 ? fifo_41_io_deqValid : 1'h0;
  assign T884 = T405 & T885;
  assign T885 = T489[3'h7:3'h7];
  assign T886 = T408 & T885;
  assign T887 = bankToPortValid_0_7;
  assign bankToPortValid_0_7 = T888;
  assign T888 = T892 ? 1'h0 : T889;
  assign T889 = T890 ? fifo_40_io_deqValid : 1'h0;
  assign T890 = T402 & T891;
  assign T891 = T497[3'h7:3'h7];
  assign T892 = T500 & T891;
  assign T893 = T894;
  assign T894 = T901 & T895;
  assign T895 = bankToPortValid_7_8;
  assign bankToPortValid_7_8 = T896;
  assign T896 = T900 ? 1'h0 : T897;
  assign T897 = T898 ? fifo_47_io_deqValid : 1'h0;
  assign T898 = T269 & T899;
  assign T899 = T368[4'h8:4'h8];
  assign T900 = T436 & T899;
  assign T901 = T908 & T902;
  assign T902 = bankToPortValid_6_8;
  assign bankToPortValid_6_8 = T903;
  assign T903 = T907 ? 1'h0 : T904;
  assign T904 = T905 ? fifo_46_io_deqValid : 1'h0;
  assign T905 = T430 & T906;
  assign T906 = T444[4'h8:4'h8];
  assign T907 = T433 & T906;
  assign T908 = T915 & T909;
  assign T909 = bankToPortValid_5_8;
  assign bankToPortValid_5_8 = T910;
  assign T910 = T914 ? 1'h0 : T911;
  assign T911 = T912 ? fifo_45_io_deqValid : 1'h0;
  assign T912 = T425 & T913;
  assign T913 = T453[4'h8:4'h8];
  assign T914 = T428 & T913;
  assign T915 = T922 & T916;
  assign T916 = bankToPortValid_4_8;
  assign bankToPortValid_4_8 = T917;
  assign T917 = T921 ? 1'h0 : T918;
  assign T918 = T919 ? fifo_44_io_deqValid : 1'h0;
  assign T919 = T420 & T920;
  assign T920 = T462[4'h8:4'h8];
  assign T921 = T423 & T920;
  assign T922 = T929 & T923;
  assign T923 = bankToPortValid_3_8;
  assign bankToPortValid_3_8 = T924;
  assign T924 = T928 ? 1'h0 : T925;
  assign T925 = T926 ? fifo_43_io_deqValid : 1'h0;
  assign T926 = T415 & T927;
  assign T927 = T471[4'h8:4'h8];
  assign T928 = T418 & T927;
  assign T929 = T936 & T930;
  assign T930 = bankToPortValid_2_8;
  assign bankToPortValid_2_8 = T931;
  assign T931 = T935 ? 1'h0 : T932;
  assign T932 = T933 ? fifo_42_io_deqValid : 1'h0;
  assign T933 = T410 & T934;
  assign T934 = T480[4'h8:4'h8];
  assign T935 = T413 & T934;
  assign T936 = T943 & T937;
  assign T937 = bankToPortValid_1_8;
  assign bankToPortValid_1_8 = T938;
  assign T938 = T942 ? 1'h0 : T939;
  assign T939 = T940 ? fifo_41_io_deqValid : 1'h0;
  assign T940 = T405 & T941;
  assign T941 = T489[4'h8:4'h8];
  assign T942 = T408 & T941;
  assign T943 = bankToPortValid_0_8;
  assign bankToPortValid_0_8 = T944;
  assign T944 = T948 ? 1'h0 : T945;
  assign T945 = T946 ? fifo_40_io_deqValid : 1'h0;
  assign T946 = T402 & T947;
  assign T947 = T497[4'h8:4'h8];
  assign T948 = T500 & T947;
  assign T949 = T950;
  assign T950 = T957 & T951;
  assign T951 = bankToPortValid_7_9;
  assign bankToPortValid_7_9 = T952;
  assign T952 = T956 ? 1'h0 : T953;
  assign T953 = T954 ? fifo_47_io_deqValid : 1'h0;
  assign T954 = T269 & T955;
  assign T955 = T368[4'h9:4'h9];
  assign T956 = T436 & T955;
  assign T957 = T964 & T958;
  assign T958 = bankToPortValid_6_9;
  assign bankToPortValid_6_9 = T959;
  assign T959 = T963 ? 1'h0 : T960;
  assign T960 = T961 ? fifo_46_io_deqValid : 1'h0;
  assign T961 = T430 & T962;
  assign T962 = T444[4'h9:4'h9];
  assign T963 = T433 & T962;
  assign T964 = T971 & T965;
  assign T965 = bankToPortValid_5_9;
  assign bankToPortValid_5_9 = T966;
  assign T966 = T970 ? 1'h0 : T967;
  assign T967 = T968 ? fifo_45_io_deqValid : 1'h0;
  assign T968 = T425 & T969;
  assign T969 = T453[4'h9:4'h9];
  assign T970 = T428 & T969;
  assign T971 = T978 & T972;
  assign T972 = bankToPortValid_4_9;
  assign bankToPortValid_4_9 = T973;
  assign T973 = T977 ? 1'h0 : T974;
  assign T974 = T975 ? fifo_44_io_deqValid : 1'h0;
  assign T975 = T420 & T976;
  assign T976 = T462[4'h9:4'h9];
  assign T977 = T423 & T976;
  assign T978 = T985 & T979;
  assign T979 = bankToPortValid_3_9;
  assign bankToPortValid_3_9 = T980;
  assign T980 = T984 ? 1'h0 : T981;
  assign T981 = T982 ? fifo_43_io_deqValid : 1'h0;
  assign T982 = T415 & T983;
  assign T983 = T471[4'h9:4'h9];
  assign T984 = T418 & T983;
  assign T985 = T992 & T986;
  assign T986 = bankToPortValid_2_9;
  assign bankToPortValid_2_9 = T987;
  assign T987 = T991 ? 1'h0 : T988;
  assign T988 = T989 ? fifo_42_io_deqValid : 1'h0;
  assign T989 = T410 & T990;
  assign T990 = T480[4'h9:4'h9];
  assign T991 = T413 & T990;
  assign T992 = T999 & T993;
  assign T993 = bankToPortValid_1_9;
  assign bankToPortValid_1_9 = T994;
  assign T994 = T998 ? 1'h0 : T995;
  assign T995 = T996 ? fifo_41_io_deqValid : 1'h0;
  assign T996 = T405 & T997;
  assign T997 = T489[4'h9:4'h9];
  assign T998 = T408 & T997;
  assign T999 = bankToPortValid_0_9;
  assign bankToPortValid_0_9 = T1000;
  assign T1000 = T1004 ? 1'h0 : T1001;
  assign T1001 = T1002 ? fifo_40_io_deqValid : 1'h0;
  assign T1002 = T402 & T1003;
  assign T1003 = T497[4'h9:4'h9];
  assign T1004 = T500 & T1003;
  assign T1005 = T1006;
  assign T1006 = T1013 & T1007;
  assign T1007 = bankToPortValid_7_10;
  assign bankToPortValid_7_10 = T1008;
  assign T1008 = T1012 ? 1'h0 : T1009;
  assign T1009 = T1010 ? fifo_47_io_deqValid : 1'h0;
  assign T1010 = T269 & T1011;
  assign T1011 = T368[4'ha:4'ha];
  assign T1012 = T436 & T1011;
  assign T1013 = T1020 & T1014;
  assign T1014 = bankToPortValid_6_10;
  assign bankToPortValid_6_10 = T1015;
  assign T1015 = T1019 ? 1'h0 : T1016;
  assign T1016 = T1017 ? fifo_46_io_deqValid : 1'h0;
  assign T1017 = T430 & T1018;
  assign T1018 = T444[4'ha:4'ha];
  assign T1019 = T433 & T1018;
  assign T1020 = T1027 & T1021;
  assign T1021 = bankToPortValid_5_10;
  assign bankToPortValid_5_10 = T1022;
  assign T1022 = T1026 ? 1'h0 : T1023;
  assign T1023 = T1024 ? fifo_45_io_deqValid : 1'h0;
  assign T1024 = T425 & T1025;
  assign T1025 = T453[4'ha:4'ha];
  assign T1026 = T428 & T1025;
  assign T1027 = T1034 & T1028;
  assign T1028 = bankToPortValid_4_10;
  assign bankToPortValid_4_10 = T1029;
  assign T1029 = T1033 ? 1'h0 : T1030;
  assign T1030 = T1031 ? fifo_44_io_deqValid : 1'h0;
  assign T1031 = T420 & T1032;
  assign T1032 = T462[4'ha:4'ha];
  assign T1033 = T423 & T1032;
  assign T1034 = T1041 & T1035;
  assign T1035 = bankToPortValid_3_10;
  assign bankToPortValid_3_10 = T1036;
  assign T1036 = T1040 ? 1'h0 : T1037;
  assign T1037 = T1038 ? fifo_43_io_deqValid : 1'h0;
  assign T1038 = T415 & T1039;
  assign T1039 = T471[4'ha:4'ha];
  assign T1040 = T418 & T1039;
  assign T1041 = T1048 & T1042;
  assign T1042 = bankToPortValid_2_10;
  assign bankToPortValid_2_10 = T1043;
  assign T1043 = T1047 ? 1'h0 : T1044;
  assign T1044 = T1045 ? fifo_42_io_deqValid : 1'h0;
  assign T1045 = T410 & T1046;
  assign T1046 = T480[4'ha:4'ha];
  assign T1047 = T413 & T1046;
  assign T1048 = T1055 & T1049;
  assign T1049 = bankToPortValid_1_10;
  assign bankToPortValid_1_10 = T1050;
  assign T1050 = T1054 ? 1'h0 : T1051;
  assign T1051 = T1052 ? fifo_41_io_deqValid : 1'h0;
  assign T1052 = T405 & T1053;
  assign T1053 = T489[4'ha:4'ha];
  assign T1054 = T408 & T1053;
  assign T1055 = bankToPortValid_0_10;
  assign bankToPortValid_0_10 = T1056;
  assign T1056 = T1060 ? 1'h0 : T1057;
  assign T1057 = T1058 ? fifo_40_io_deqValid : 1'h0;
  assign T1058 = T402 & T1059;
  assign T1059 = T497[4'ha:4'ha];
  assign T1060 = T500 & T1059;
  assign T1061 = T1062;
  assign T1062 = T1069 & T1063;
  assign T1063 = bankToPortValid_7_11;
  assign bankToPortValid_7_11 = T1064;
  assign T1064 = T1068 ? 1'h0 : T1065;
  assign T1065 = T1066 ? fifo_47_io_deqValid : 1'h0;
  assign T1066 = T269 & T1067;
  assign T1067 = T368[4'hb:4'hb];
  assign T1068 = T436 & T1067;
  assign T1069 = T1076 & T1070;
  assign T1070 = bankToPortValid_6_11;
  assign bankToPortValid_6_11 = T1071;
  assign T1071 = T1075 ? 1'h0 : T1072;
  assign T1072 = T1073 ? fifo_46_io_deqValid : 1'h0;
  assign T1073 = T430 & T1074;
  assign T1074 = T444[4'hb:4'hb];
  assign T1075 = T433 & T1074;
  assign T1076 = T1083 & T1077;
  assign T1077 = bankToPortValid_5_11;
  assign bankToPortValid_5_11 = T1078;
  assign T1078 = T1082 ? 1'h0 : T1079;
  assign T1079 = T1080 ? fifo_45_io_deqValid : 1'h0;
  assign T1080 = T425 & T1081;
  assign T1081 = T453[4'hb:4'hb];
  assign T1082 = T428 & T1081;
  assign T1083 = T1090 & T1084;
  assign T1084 = bankToPortValid_4_11;
  assign bankToPortValid_4_11 = T1085;
  assign T1085 = T1089 ? 1'h0 : T1086;
  assign T1086 = T1087 ? fifo_44_io_deqValid : 1'h0;
  assign T1087 = T420 & T1088;
  assign T1088 = T462[4'hb:4'hb];
  assign T1089 = T423 & T1088;
  assign T1090 = T1097 & T1091;
  assign T1091 = bankToPortValid_3_11;
  assign bankToPortValid_3_11 = T1092;
  assign T1092 = T1096 ? 1'h0 : T1093;
  assign T1093 = T1094 ? fifo_43_io_deqValid : 1'h0;
  assign T1094 = T415 & T1095;
  assign T1095 = T471[4'hb:4'hb];
  assign T1096 = T418 & T1095;
  assign T1097 = T1104 & T1098;
  assign T1098 = bankToPortValid_2_11;
  assign bankToPortValid_2_11 = T1099;
  assign T1099 = T1103 ? 1'h0 : T1100;
  assign T1100 = T1101 ? fifo_42_io_deqValid : 1'h0;
  assign T1101 = T410 & T1102;
  assign T1102 = T480[4'hb:4'hb];
  assign T1103 = T413 & T1102;
  assign T1104 = T1111 & T1105;
  assign T1105 = bankToPortValid_1_11;
  assign bankToPortValid_1_11 = T1106;
  assign T1106 = T1110 ? 1'h0 : T1107;
  assign T1107 = T1108 ? fifo_41_io_deqValid : 1'h0;
  assign T1108 = T405 & T1109;
  assign T1109 = T489[4'hb:4'hb];
  assign T1110 = T408 & T1109;
  assign T1111 = bankToPortValid_0_11;
  assign bankToPortValid_0_11 = T1112;
  assign T1112 = T1116 ? 1'h0 : T1113;
  assign T1113 = T1114 ? fifo_40_io_deqValid : 1'h0;
  assign T1114 = T402 & T1115;
  assign T1115 = T497[4'hb:4'hb];
  assign T1116 = T500 & T1115;
  assign T1117 = T1118;
  assign T1118 = T1125 & T1119;
  assign T1119 = bankToPortValid_7_12;
  assign bankToPortValid_7_12 = T1120;
  assign T1120 = T1124 ? 1'h0 : T1121;
  assign T1121 = T1122 ? fifo_47_io_deqValid : 1'h0;
  assign T1122 = T269 & T1123;
  assign T1123 = T368[4'hc:4'hc];
  assign T1124 = T436 & T1123;
  assign T1125 = T1132 & T1126;
  assign T1126 = bankToPortValid_6_12;
  assign bankToPortValid_6_12 = T1127;
  assign T1127 = T1131 ? 1'h0 : T1128;
  assign T1128 = T1129 ? fifo_46_io_deqValid : 1'h0;
  assign T1129 = T430 & T1130;
  assign T1130 = T444[4'hc:4'hc];
  assign T1131 = T433 & T1130;
  assign T1132 = T1139 & T1133;
  assign T1133 = bankToPortValid_5_12;
  assign bankToPortValid_5_12 = T1134;
  assign T1134 = T1138 ? 1'h0 : T1135;
  assign T1135 = T1136 ? fifo_45_io_deqValid : 1'h0;
  assign T1136 = T425 & T1137;
  assign T1137 = T453[4'hc:4'hc];
  assign T1138 = T428 & T1137;
  assign T1139 = T1146 & T1140;
  assign T1140 = bankToPortValid_4_12;
  assign bankToPortValid_4_12 = T1141;
  assign T1141 = T1145 ? 1'h0 : T1142;
  assign T1142 = T1143 ? fifo_44_io_deqValid : 1'h0;
  assign T1143 = T420 & T1144;
  assign T1144 = T462[4'hc:4'hc];
  assign T1145 = T423 & T1144;
  assign T1146 = T1153 & T1147;
  assign T1147 = bankToPortValid_3_12;
  assign bankToPortValid_3_12 = T1148;
  assign T1148 = T1152 ? 1'h0 : T1149;
  assign T1149 = T1150 ? fifo_43_io_deqValid : 1'h0;
  assign T1150 = T415 & T1151;
  assign T1151 = T471[4'hc:4'hc];
  assign T1152 = T418 & T1151;
  assign T1153 = T1160 & T1154;
  assign T1154 = bankToPortValid_2_12;
  assign bankToPortValid_2_12 = T1155;
  assign T1155 = T1159 ? 1'h0 : T1156;
  assign T1156 = T1157 ? fifo_42_io_deqValid : 1'h0;
  assign T1157 = T410 & T1158;
  assign T1158 = T480[4'hc:4'hc];
  assign T1159 = T413 & T1158;
  assign T1160 = T1167 & T1161;
  assign T1161 = bankToPortValid_1_12;
  assign bankToPortValid_1_12 = T1162;
  assign T1162 = T1166 ? 1'h0 : T1163;
  assign T1163 = T1164 ? fifo_41_io_deqValid : 1'h0;
  assign T1164 = T405 & T1165;
  assign T1165 = T489[4'hc:4'hc];
  assign T1166 = T408 & T1165;
  assign T1167 = bankToPortValid_0_12;
  assign bankToPortValid_0_12 = T1168;
  assign T1168 = T1172 ? 1'h0 : T1169;
  assign T1169 = T1170 ? fifo_40_io_deqValid : 1'h0;
  assign T1170 = T402 & T1171;
  assign T1171 = T497[4'hc:4'hc];
  assign T1172 = T500 & T1171;
  assign T1173 = T1174;
  assign T1174 = T1181 & T1175;
  assign T1175 = bankToPortValid_7_13;
  assign bankToPortValid_7_13 = T1176;
  assign T1176 = T1180 ? 1'h0 : T1177;
  assign T1177 = T1178 ? fifo_47_io_deqValid : 1'h0;
  assign T1178 = T269 & T1179;
  assign T1179 = T368[4'hd:4'hd];
  assign T1180 = T436 & T1179;
  assign T1181 = T1188 & T1182;
  assign T1182 = bankToPortValid_6_13;
  assign bankToPortValid_6_13 = T1183;
  assign T1183 = T1187 ? 1'h0 : T1184;
  assign T1184 = T1185 ? fifo_46_io_deqValid : 1'h0;
  assign T1185 = T430 & T1186;
  assign T1186 = T444[4'hd:4'hd];
  assign T1187 = T433 & T1186;
  assign T1188 = T1195 & T1189;
  assign T1189 = bankToPortValid_5_13;
  assign bankToPortValid_5_13 = T1190;
  assign T1190 = T1194 ? 1'h0 : T1191;
  assign T1191 = T1192 ? fifo_45_io_deqValid : 1'h0;
  assign T1192 = T425 & T1193;
  assign T1193 = T453[4'hd:4'hd];
  assign T1194 = T428 & T1193;
  assign T1195 = T1202 & T1196;
  assign T1196 = bankToPortValid_4_13;
  assign bankToPortValid_4_13 = T1197;
  assign T1197 = T1201 ? 1'h0 : T1198;
  assign T1198 = T1199 ? fifo_44_io_deqValid : 1'h0;
  assign T1199 = T420 & T1200;
  assign T1200 = T462[4'hd:4'hd];
  assign T1201 = T423 & T1200;
  assign T1202 = T1209 & T1203;
  assign T1203 = bankToPortValid_3_13;
  assign bankToPortValid_3_13 = T1204;
  assign T1204 = T1208 ? 1'h0 : T1205;
  assign T1205 = T1206 ? fifo_43_io_deqValid : 1'h0;
  assign T1206 = T415 & T1207;
  assign T1207 = T471[4'hd:4'hd];
  assign T1208 = T418 & T1207;
  assign T1209 = T1216 & T1210;
  assign T1210 = bankToPortValid_2_13;
  assign bankToPortValid_2_13 = T1211;
  assign T1211 = T1215 ? 1'h0 : T1212;
  assign T1212 = T1213 ? fifo_42_io_deqValid : 1'h0;
  assign T1213 = T410 & T1214;
  assign T1214 = T480[4'hd:4'hd];
  assign T1215 = T413 & T1214;
  assign T1216 = T1223 & T1217;
  assign T1217 = bankToPortValid_1_13;
  assign bankToPortValid_1_13 = T1218;
  assign T1218 = T1222 ? 1'h0 : T1219;
  assign T1219 = T1220 ? fifo_41_io_deqValid : 1'h0;
  assign T1220 = T405 & T1221;
  assign T1221 = T489[4'hd:4'hd];
  assign T1222 = T408 & T1221;
  assign T1223 = bankToPortValid_0_13;
  assign bankToPortValid_0_13 = T1224;
  assign T1224 = T1228 ? 1'h0 : T1225;
  assign T1225 = T1226 ? fifo_40_io_deqValid : 1'h0;
  assign T1226 = T402 & T1227;
  assign T1227 = T497[4'hd:4'hd];
  assign T1228 = T500 & T1227;
  assign T1229 = T1230;
  assign T1230 = T1237 & T1231;
  assign T1231 = bankToPortValid_7_14;
  assign bankToPortValid_7_14 = T1232;
  assign T1232 = T1236 ? 1'h0 : T1233;
  assign T1233 = T1234 ? fifo_47_io_deqValid : 1'h0;
  assign T1234 = T269 & T1235;
  assign T1235 = T368[4'he:4'he];
  assign T1236 = T436 & T1235;
  assign T1237 = T1244 & T1238;
  assign T1238 = bankToPortValid_6_14;
  assign bankToPortValid_6_14 = T1239;
  assign T1239 = T1243 ? 1'h0 : T1240;
  assign T1240 = T1241 ? fifo_46_io_deqValid : 1'h0;
  assign T1241 = T430 & T1242;
  assign T1242 = T444[4'he:4'he];
  assign T1243 = T433 & T1242;
  assign T1244 = T1251 & T1245;
  assign T1245 = bankToPortValid_5_14;
  assign bankToPortValid_5_14 = T1246;
  assign T1246 = T1250 ? 1'h0 : T1247;
  assign T1247 = T1248 ? fifo_45_io_deqValid : 1'h0;
  assign T1248 = T425 & T1249;
  assign T1249 = T453[4'he:4'he];
  assign T1250 = T428 & T1249;
  assign T1251 = T1258 & T1252;
  assign T1252 = bankToPortValid_4_14;
  assign bankToPortValid_4_14 = T1253;
  assign T1253 = T1257 ? 1'h0 : T1254;
  assign T1254 = T1255 ? fifo_44_io_deqValid : 1'h0;
  assign T1255 = T420 & T1256;
  assign T1256 = T462[4'he:4'he];
  assign T1257 = T423 & T1256;
  assign T1258 = T1265 & T1259;
  assign T1259 = bankToPortValid_3_14;
  assign bankToPortValid_3_14 = T1260;
  assign T1260 = T1264 ? 1'h0 : T1261;
  assign T1261 = T1262 ? fifo_43_io_deqValid : 1'h0;
  assign T1262 = T415 & T1263;
  assign T1263 = T471[4'he:4'he];
  assign T1264 = T418 & T1263;
  assign T1265 = T1272 & T1266;
  assign T1266 = bankToPortValid_2_14;
  assign bankToPortValid_2_14 = T1267;
  assign T1267 = T1271 ? 1'h0 : T1268;
  assign T1268 = T1269 ? fifo_42_io_deqValid : 1'h0;
  assign T1269 = T410 & T1270;
  assign T1270 = T480[4'he:4'he];
  assign T1271 = T413 & T1270;
  assign T1272 = T1279 & T1273;
  assign T1273 = bankToPortValid_1_14;
  assign bankToPortValid_1_14 = T1274;
  assign T1274 = T1278 ? 1'h0 : T1275;
  assign T1275 = T1276 ? fifo_41_io_deqValid : 1'h0;
  assign T1276 = T405 & T1277;
  assign T1277 = T489[4'he:4'he];
  assign T1278 = T408 & T1277;
  assign T1279 = bankToPortValid_0_14;
  assign bankToPortValid_0_14 = T1280;
  assign T1280 = T1284 ? 1'h0 : T1281;
  assign T1281 = T1282 ? fifo_40_io_deqValid : 1'h0;
  assign T1282 = T402 & T1283;
  assign T1283 = T497[4'he:4'he];
  assign T1284 = T500 & T1283;
  assign T1285 = T1286;
  assign T1286 = T1293 & T1287;
  assign T1287 = bankToPortValid_7_15;
  assign bankToPortValid_7_15 = T1288;
  assign T1288 = T1292 ? 1'h0 : T1289;
  assign T1289 = T1290 ? fifo_47_io_deqValid : 1'h0;
  assign T1290 = T269 & T1291;
  assign T1291 = T368[4'hf:4'hf];
  assign T1292 = T436 & T1291;
  assign T1293 = T1300 & T1294;
  assign T1294 = bankToPortValid_6_15;
  assign bankToPortValid_6_15 = T1295;
  assign T1295 = T1299 ? 1'h0 : T1296;
  assign T1296 = T1297 ? fifo_46_io_deqValid : 1'h0;
  assign T1297 = T430 & T1298;
  assign T1298 = T444[4'hf:4'hf];
  assign T1299 = T433 & T1298;
  assign T1300 = T1307 & T1301;
  assign T1301 = bankToPortValid_5_15;
  assign bankToPortValid_5_15 = T1302;
  assign T1302 = T1306 ? 1'h0 : T1303;
  assign T1303 = T1304 ? fifo_45_io_deqValid : 1'h0;
  assign T1304 = T425 & T1305;
  assign T1305 = T453[4'hf:4'hf];
  assign T1306 = T428 & T1305;
  assign T1307 = T1314 & T1308;
  assign T1308 = bankToPortValid_4_15;
  assign bankToPortValid_4_15 = T1309;
  assign T1309 = T1313 ? 1'h0 : T1310;
  assign T1310 = T1311 ? fifo_44_io_deqValid : 1'h0;
  assign T1311 = T420 & T1312;
  assign T1312 = T462[4'hf:4'hf];
  assign T1313 = T423 & T1312;
  assign T1314 = T1321 & T1315;
  assign T1315 = bankToPortValid_3_15;
  assign bankToPortValid_3_15 = T1316;
  assign T1316 = T1320 ? 1'h0 : T1317;
  assign T1317 = T1318 ? fifo_43_io_deqValid : 1'h0;
  assign T1318 = T415 & T1319;
  assign T1319 = T471[4'hf:4'hf];
  assign T1320 = T418 & T1319;
  assign T1321 = T1328 & T1322;
  assign T1322 = bankToPortValid_2_15;
  assign bankToPortValid_2_15 = T1323;
  assign T1323 = T1327 ? 1'h0 : T1324;
  assign T1324 = T1325 ? fifo_42_io_deqValid : 1'h0;
  assign T1325 = T410 & T1326;
  assign T1326 = T480[4'hf:4'hf];
  assign T1327 = T413 & T1326;
  assign T1328 = T1335 & T1329;
  assign T1329 = bankToPortValid_1_15;
  assign bankToPortValid_1_15 = T1330;
  assign T1330 = T1334 ? 1'h0 : T1331;
  assign T1331 = T1332 ? fifo_41_io_deqValid : 1'h0;
  assign T1332 = T405 & T1333;
  assign T1333 = T489[4'hf:4'hf];
  assign T1334 = T408 & T1333;
  assign T1335 = bankToPortValid_0_15;
  assign bankToPortValid_0_15 = T1336;
  assign T1336 = T1340 ? 1'h0 : T1337;
  assign T1337 = T1338 ? fifo_40_io_deqValid : 1'h0;
  assign T1338 = T402 & T1339;
  assign T1339 = T497[4'hf:4'hf];
  assign T1340 = T500 & T1339;
  assign T1341 = T1342;
  assign T1342 = T1349 & T1343;
  assign T1343 = bankToPortValid_7_16;
  assign bankToPortValid_7_16 = T1344;
  assign T1344 = T1348 ? 1'h0 : T1345;
  assign T1345 = T1346 ? fifo_47_io_deqValid : 1'h0;
  assign T1346 = T269 & T1347;
  assign T1347 = T368[5'h10:5'h10];
  assign T1348 = T436 & T1347;
  assign T1349 = T1356 & T1350;
  assign T1350 = bankToPortValid_6_16;
  assign bankToPortValid_6_16 = T1351;
  assign T1351 = T1355 ? 1'h0 : T1352;
  assign T1352 = T1353 ? fifo_46_io_deqValid : 1'h0;
  assign T1353 = T430 & T1354;
  assign T1354 = T444[5'h10:5'h10];
  assign T1355 = T433 & T1354;
  assign T1356 = T1363 & T1357;
  assign T1357 = bankToPortValid_5_16;
  assign bankToPortValid_5_16 = T1358;
  assign T1358 = T1362 ? 1'h0 : T1359;
  assign T1359 = T1360 ? fifo_45_io_deqValid : 1'h0;
  assign T1360 = T425 & T1361;
  assign T1361 = T453[5'h10:5'h10];
  assign T1362 = T428 & T1361;
  assign T1363 = T1370 & T1364;
  assign T1364 = bankToPortValid_4_16;
  assign bankToPortValid_4_16 = T1365;
  assign T1365 = T1369 ? 1'h0 : T1366;
  assign T1366 = T1367 ? fifo_44_io_deqValid : 1'h0;
  assign T1367 = T420 & T1368;
  assign T1368 = T462[5'h10:5'h10];
  assign T1369 = T423 & T1368;
  assign T1370 = T1377 & T1371;
  assign T1371 = bankToPortValid_3_16;
  assign bankToPortValid_3_16 = T1372;
  assign T1372 = T1376 ? 1'h0 : T1373;
  assign T1373 = T1374 ? fifo_43_io_deqValid : 1'h0;
  assign T1374 = T415 & T1375;
  assign T1375 = T471[5'h10:5'h10];
  assign T1376 = T418 & T1375;
  assign T1377 = T1384 & T1378;
  assign T1378 = bankToPortValid_2_16;
  assign bankToPortValid_2_16 = T1379;
  assign T1379 = T1383 ? 1'h0 : T1380;
  assign T1380 = T1381 ? fifo_42_io_deqValid : 1'h0;
  assign T1381 = T410 & T1382;
  assign T1382 = T480[5'h10:5'h10];
  assign T1383 = T413 & T1382;
  assign T1384 = T1391 & T1385;
  assign T1385 = bankToPortValid_1_16;
  assign bankToPortValid_1_16 = T1386;
  assign T1386 = T1390 ? 1'h0 : T1387;
  assign T1387 = T1388 ? fifo_41_io_deqValid : 1'h0;
  assign T1388 = T405 & T1389;
  assign T1389 = T489[5'h10:5'h10];
  assign T1390 = T408 & T1389;
  assign T1391 = bankToPortValid_0_16;
  assign bankToPortValid_0_16 = T1392;
  assign T1392 = T1396 ? 1'h0 : T1393;
  assign T1393 = T1394 ? fifo_40_io_deqValid : 1'h0;
  assign T1394 = T402 & T1395;
  assign T1395 = T497[5'h10:5'h10];
  assign T1396 = T500 & T1395;
  assign T1397 = T1398;
  assign T1398 = T1405 & T1399;
  assign T1399 = bankToPortValid_7_17;
  assign bankToPortValid_7_17 = T1400;
  assign T1400 = T1404 ? 1'h0 : T1401;
  assign T1401 = T1402 ? fifo_47_io_deqValid : 1'h0;
  assign T1402 = T269 & T1403;
  assign T1403 = T368[5'h11:5'h11];
  assign T1404 = T436 & T1403;
  assign T1405 = T1412 & T1406;
  assign T1406 = bankToPortValid_6_17;
  assign bankToPortValid_6_17 = T1407;
  assign T1407 = T1411 ? 1'h0 : T1408;
  assign T1408 = T1409 ? fifo_46_io_deqValid : 1'h0;
  assign T1409 = T430 & T1410;
  assign T1410 = T444[5'h11:5'h11];
  assign T1411 = T433 & T1410;
  assign T1412 = T1419 & T1413;
  assign T1413 = bankToPortValid_5_17;
  assign bankToPortValid_5_17 = T1414;
  assign T1414 = T1418 ? 1'h0 : T1415;
  assign T1415 = T1416 ? fifo_45_io_deqValid : 1'h0;
  assign T1416 = T425 & T1417;
  assign T1417 = T453[5'h11:5'h11];
  assign T1418 = T428 & T1417;
  assign T1419 = T1426 & T1420;
  assign T1420 = bankToPortValid_4_17;
  assign bankToPortValid_4_17 = T1421;
  assign T1421 = T1425 ? 1'h0 : T1422;
  assign T1422 = T1423 ? fifo_44_io_deqValid : 1'h0;
  assign T1423 = T420 & T1424;
  assign T1424 = T462[5'h11:5'h11];
  assign T1425 = T423 & T1424;
  assign T1426 = T1433 & T1427;
  assign T1427 = bankToPortValid_3_17;
  assign bankToPortValid_3_17 = T1428;
  assign T1428 = T1432 ? 1'h0 : T1429;
  assign T1429 = T1430 ? fifo_43_io_deqValid : 1'h0;
  assign T1430 = T415 & T1431;
  assign T1431 = T471[5'h11:5'h11];
  assign T1432 = T418 & T1431;
  assign T1433 = T1440 & T1434;
  assign T1434 = bankToPortValid_2_17;
  assign bankToPortValid_2_17 = T1435;
  assign T1435 = T1439 ? 1'h0 : T1436;
  assign T1436 = T1437 ? fifo_42_io_deqValid : 1'h0;
  assign T1437 = T410 & T1438;
  assign T1438 = T480[5'h11:5'h11];
  assign T1439 = T413 & T1438;
  assign T1440 = T1447 & T1441;
  assign T1441 = bankToPortValid_1_17;
  assign bankToPortValid_1_17 = T1442;
  assign T1442 = T1446 ? 1'h0 : T1443;
  assign T1443 = T1444 ? fifo_41_io_deqValid : 1'h0;
  assign T1444 = T405 & T1445;
  assign T1445 = T489[5'h11:5'h11];
  assign T1446 = T408 & T1445;
  assign T1447 = bankToPortValid_0_17;
  assign bankToPortValid_0_17 = T1448;
  assign T1448 = T1452 ? 1'h0 : T1449;
  assign T1449 = T1450 ? fifo_40_io_deqValid : 1'h0;
  assign T1450 = T402 & T1451;
  assign T1451 = T497[5'h11:5'h11];
  assign T1452 = T500 & T1451;
  assign T1453 = T1454;
  assign T1454 = T1461 & T1455;
  assign T1455 = bankToPortValid_7_18;
  assign bankToPortValid_7_18 = T1456;
  assign T1456 = T1460 ? 1'h0 : T1457;
  assign T1457 = T1458 ? fifo_47_io_deqValid : 1'h0;
  assign T1458 = T269 & T1459;
  assign T1459 = T368[5'h12:5'h12];
  assign T1460 = T436 & T1459;
  assign T1461 = T1468 & T1462;
  assign T1462 = bankToPortValid_6_18;
  assign bankToPortValid_6_18 = T1463;
  assign T1463 = T1467 ? 1'h0 : T1464;
  assign T1464 = T1465 ? fifo_46_io_deqValid : 1'h0;
  assign T1465 = T430 & T1466;
  assign T1466 = T444[5'h12:5'h12];
  assign T1467 = T433 & T1466;
  assign T1468 = T1475 & T1469;
  assign T1469 = bankToPortValid_5_18;
  assign bankToPortValid_5_18 = T1470;
  assign T1470 = T1474 ? 1'h0 : T1471;
  assign T1471 = T1472 ? fifo_45_io_deqValid : 1'h0;
  assign T1472 = T425 & T1473;
  assign T1473 = T453[5'h12:5'h12];
  assign T1474 = T428 & T1473;
  assign T1475 = T1482 & T1476;
  assign T1476 = bankToPortValid_4_18;
  assign bankToPortValid_4_18 = T1477;
  assign T1477 = T1481 ? 1'h0 : T1478;
  assign T1478 = T1479 ? fifo_44_io_deqValid : 1'h0;
  assign T1479 = T420 & T1480;
  assign T1480 = T462[5'h12:5'h12];
  assign T1481 = T423 & T1480;
  assign T1482 = T1489 & T1483;
  assign T1483 = bankToPortValid_3_18;
  assign bankToPortValid_3_18 = T1484;
  assign T1484 = T1488 ? 1'h0 : T1485;
  assign T1485 = T1486 ? fifo_43_io_deqValid : 1'h0;
  assign T1486 = T415 & T1487;
  assign T1487 = T471[5'h12:5'h12];
  assign T1488 = T418 & T1487;
  assign T1489 = T1496 & T1490;
  assign T1490 = bankToPortValid_2_18;
  assign bankToPortValid_2_18 = T1491;
  assign T1491 = T1495 ? 1'h0 : T1492;
  assign T1492 = T1493 ? fifo_42_io_deqValid : 1'h0;
  assign T1493 = T410 & T1494;
  assign T1494 = T480[5'h12:5'h12];
  assign T1495 = T413 & T1494;
  assign T1496 = T1503 & T1497;
  assign T1497 = bankToPortValid_1_18;
  assign bankToPortValid_1_18 = T1498;
  assign T1498 = T1502 ? 1'h0 : T1499;
  assign T1499 = T1500 ? fifo_41_io_deqValid : 1'h0;
  assign T1500 = T405 & T1501;
  assign T1501 = T489[5'h12:5'h12];
  assign T1502 = T408 & T1501;
  assign T1503 = bankToPortValid_0_18;
  assign bankToPortValid_0_18 = T1504;
  assign T1504 = T1508 ? 1'h0 : T1505;
  assign T1505 = T1506 ? fifo_40_io_deqValid : 1'h0;
  assign T1506 = T402 & T1507;
  assign T1507 = T497[5'h12:5'h12];
  assign T1508 = T500 & T1507;
  assign T3128 = reset ? 1'h0 : T336;
  assign T336 = fabInSeqMemConfig_io_rst ? 1'h0 : T337;
  assign T337 = T67 ? T359 : T338;
  assign T338 = T78 ? T357 : T339;
  assign T339 = T89 ? T355 : T340;
  assign T340 = T100 ? T353 : T341;
  assign T341 = T111 ? T351 : T342;
  assign T342 = T122 ? T349 : T343;
  assign T343 = T133 ? T347 : T344;
  assign T344 = T143 ? T345 : seqLevelDoneReg1;
  assign T345 = ~ T346;
  assign T346 = nextSeq[7'h58:7'h58];
  assign T347 = ~ T348;
  assign T348 = nextSeq[7'h58:7'h58];
  assign T349 = ~ T350;
  assign T350 = nextSeq[7'h58:7'h58];
  assign T351 = ~ T352;
  assign T352 = nextSeq[7'h58:7'h58];
  assign T353 = ~ T354;
  assign T354 = nextSeq[7'h58:7'h58];
  assign T355 = ~ T356;
  assign T356 = nextSeq[7'h58:7'h58];
  assign T357 = ~ T358;
  assign T358 = nextSeq[7'h58:7'h58];
  assign T359 = ~ T360;
  assign T360 = nextSeq[7'h58:7'h58];
  assign T1509 = T1510;
  assign T1510 = T1517 & T1511;
  assign T1511 = bankToPortValid_7_19;
  assign bankToPortValid_7_19 = T1512;
  assign T1512 = T1516 ? 1'h0 : T1513;
  assign T1513 = T1514 ? fifo_47_io_deqValid : 1'h0;
  assign T1514 = T269 & T1515;
  assign T1515 = T368[5'h13:5'h13];
  assign T1516 = T436 & T1515;
  assign T1517 = T1524 & T1518;
  assign T1518 = bankToPortValid_6_19;
  assign bankToPortValid_6_19 = T1519;
  assign T1519 = T1523 ? 1'h0 : T1520;
  assign T1520 = T1521 ? fifo_46_io_deqValid : 1'h0;
  assign T1521 = T430 & T1522;
  assign T1522 = T444[5'h13:5'h13];
  assign T1523 = T433 & T1522;
  assign T1524 = T1531 & T1525;
  assign T1525 = bankToPortValid_5_19;
  assign bankToPortValid_5_19 = T1526;
  assign T1526 = T1530 ? 1'h0 : T1527;
  assign T1527 = T1528 ? fifo_45_io_deqValid : 1'h0;
  assign T1528 = T425 & T1529;
  assign T1529 = T453[5'h13:5'h13];
  assign T1530 = T428 & T1529;
  assign T1531 = T1538 & T1532;
  assign T1532 = bankToPortValid_4_19;
  assign bankToPortValid_4_19 = T1533;
  assign T1533 = T1537 ? 1'h0 : T1534;
  assign T1534 = T1535 ? fifo_44_io_deqValid : 1'h0;
  assign T1535 = T420 & T1536;
  assign T1536 = T462[5'h13:5'h13];
  assign T1537 = T423 & T1536;
  assign T1538 = T1545 & T1539;
  assign T1539 = bankToPortValid_3_19;
  assign bankToPortValid_3_19 = T1540;
  assign T1540 = T1544 ? 1'h0 : T1541;
  assign T1541 = T1542 ? fifo_43_io_deqValid : 1'h0;
  assign T1542 = T415 & T1543;
  assign T1543 = T471[5'h13:5'h13];
  assign T1544 = T418 & T1543;
  assign T1545 = T1552 & T1546;
  assign T1546 = bankToPortValid_2_19;
  assign bankToPortValid_2_19 = T1547;
  assign T1547 = T1551 ? 1'h0 : T1548;
  assign T1548 = T1549 ? fifo_42_io_deqValid : 1'h0;
  assign T1549 = T410 & T1550;
  assign T1550 = T480[5'h13:5'h13];
  assign T1551 = T413 & T1550;
  assign T1552 = T1559 & T1553;
  assign T1553 = bankToPortValid_1_19;
  assign bankToPortValid_1_19 = T1554;
  assign T1554 = T1558 ? 1'h0 : T1555;
  assign T1555 = T1556 ? fifo_41_io_deqValid : 1'h0;
  assign T1556 = T405 & T1557;
  assign T1557 = T489[5'h13:5'h13];
  assign T1558 = T408 & T1557;
  assign T1559 = bankToPortValid_0_19;
  assign bankToPortValid_0_19 = T1560;
  assign T1560 = T1564 ? 1'h0 : T1561;
  assign T1561 = T1562 ? fifo_40_io_deqValid : 1'h0;
  assign T1562 = T402 & T1563;
  assign T1563 = T497[5'h13:5'h13];
  assign T1564 = T500 & T1563;
  assign T1565 = seqLevelDoneReg2 & T1566;
  assign T1566 = rdy ^ 1'h1;
  assign T1567 = seqLevelDoneReg2 ^ 1'h1;
  assign T1568 = ~ seqLevelDoneReg2;
  assign T1569 = T267 ? readValuelocStrg : readValuelocStrg;
  assign readValuelocStrg = T3129;
  assign T3129 = T1570[5'h1f:1'h0];
  assign T1570 = T266 ? localStorage_io_outData_7 : T1571;
  assign T1571 = T267 ? localStorage_io_outData_7 : T1572;
  assign T1572 = T265 ? localStorage_io_outData_6 : T1573;
  assign T1573 = T264 ? localStorage_io_outData_6 : T1574;
  assign T1574 = T263 ? localStorage_io_outData_5 : T1575;
  assign T1575 = T262 ? localStorage_io_outData_5 : T1576;
  assign T1576 = T261 ? localStorage_io_outData_4 : T1577;
  assign T1577 = T260 ? localStorage_io_outData_4 : T1578;
  assign T1578 = T259 ? localStorage_io_outData_3 : T1579;
  assign T1579 = T258 ? localStorage_io_outData_3 : T1580;
  assign T1580 = T257 ? localStorage_io_outData_2 : T1581;
  assign T1581 = T256 ? localStorage_io_outData_2 : T1582;
  assign T1582 = T255 ? localStorage_io_outData_1 : T1583;
  assign T1583 = T254 ? localStorage_io_outData_1 : T1584;
  assign T1584 = T17 ? localStorage_io_outData_0 : localStorage_io_outData_0;
  assign T1585 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1586 = T264 ? isReadValid : 1'h0;
  assign T1587 = T430 ? 1'h1 : 1'h0;
  assign T1588 = T264 ? readValuelocStrg : readValuelocStrg;
  assign T1589 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1590 = T262 ? isReadValid : 1'h0;
  assign T1591 = T425 ? 1'h1 : 1'h0;
  assign T1592 = T262 ? readValuelocStrg : readValuelocStrg;
  assign T1593 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1594 = T260 ? isReadValid : 1'h0;
  assign T1595 = T420 ? 1'h1 : 1'h0;
  assign T1596 = T260 ? readValuelocStrg : readValuelocStrg;
  assign T1597 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1598 = T258 ? isReadValid : 1'h0;
  assign T1599 = T415 ? 1'h1 : 1'h0;
  assign T1600 = T258 ? readValuelocStrg : readValuelocStrg;
  assign T1601 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1602 = T256 ? isReadValid : 1'h0;
  assign T1603 = T410 ? 1'h1 : 1'h0;
  assign T1604 = T256 ? readValuelocStrg : readValuelocStrg;
  assign T1605 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1606 = T254 ? isReadValid : 1'h0;
  assign T1607 = T405 ? 1'h1 : 1'h0;
  assign T1608 = T254 ? readValuelocStrg : readValuelocStrg;
  assign T1609 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1610 = T17 ? isReadValid : 1'h0;
  assign T1611 = T402 ? 1'h1 : 1'h0;
  assign T1612 = T17 ? readValuelocStrg : readValuelocStrg;
  assign T1613 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1614 = T1615 ? 1'h1 : 1'h0;
  assign T1615 = T1509 & fifo_39_io_enqRdy;
  assign T1616 = seqLevelDoneReg2 ? fifo_19_io_enqRdy : 1'h0;
  assign T1617 = T1615 ? T1618 : T1618;
  assign T1618 = T1619;
  assign T1619 = T1708 ? 32'h0 : T1620;
  assign T1620 = T1509 ? T1621 : 32'h0;
  assign T1621 = T1645 | T1622;
  assign T1622 = bankToPort_7_19;
  assign bankToPort_7_19 = T1623;
  assign T1623 = T1644 ? readValueBankFifo : T1624;
  assign T1624 = T1625 ? readValueBankFifo : 32'h0;
  assign T1625 = T269 & T1626;
  assign T1626 = T1627[5'h13:5'h13];
  assign T1627 = 1'h1 << T1628;
  assign T1628 = T3130;
  assign T3130 = {2'h0, portId};
  assign readValueBankFifo = T1629;
  assign T1629 = T436 ? fifo_47_io_deqData : T1630;
  assign T1630 = T269 ? fifo_47_io_deqData : T1631;
  assign T1631 = T433 ? fifo_46_io_deqData : T1632;
  assign T1632 = T430 ? fifo_46_io_deqData : T1633;
  assign T1633 = T428 ? fifo_45_io_deqData : T1634;
  assign T1634 = T425 ? fifo_45_io_deqData : T1635;
  assign T1635 = T423 ? fifo_44_io_deqData : T1636;
  assign T1636 = T420 ? fifo_44_io_deqData : T1637;
  assign T1637 = T418 ? fifo_43_io_deqData : T1638;
  assign T1638 = T415 ? fifo_43_io_deqData : T1639;
  assign T1639 = T413 ? fifo_42_io_deqData : T1640;
  assign T1640 = T410 ? fifo_42_io_deqData : T1641;
  assign T1641 = T408 ? fifo_41_io_deqData : T1642;
  assign T1642 = T405 ? fifo_41_io_deqData : T1643;
  assign T1643 = T402 ? fifo_40_io_deqData : fifo_40_io_deqData;
  assign T1644 = T436 & T1626;
  assign T1645 = T1654 | T1646;
  assign T1646 = bankToPort_6_19;
  assign bankToPort_6_19 = T1647;
  assign T1647 = T1653 ? readValueBankFifo : T1648;
  assign T1648 = T1649 ? readValueBankFifo : 32'h0;
  assign T1649 = T430 & T1650;
  assign T1650 = T1651[5'h13:5'h13];
  assign T1651 = 1'h1 << T1652;
  assign T1652 = T3131;
  assign T3131 = {2'h0, portId};
  assign T1653 = T433 & T1650;
  assign T1654 = T1663 | T1655;
  assign T1655 = bankToPort_5_19;
  assign bankToPort_5_19 = T1656;
  assign T1656 = T1662 ? readValueBankFifo : T1657;
  assign T1657 = T1658 ? readValueBankFifo : 32'h0;
  assign T1658 = T425 & T1659;
  assign T1659 = T1660[5'h13:5'h13];
  assign T1660 = 1'h1 << T1661;
  assign T1661 = T3132;
  assign T3132 = {2'h0, portId};
  assign T1662 = T428 & T1659;
  assign T1663 = T1672 | T1664;
  assign T1664 = bankToPort_4_19;
  assign bankToPort_4_19 = T1665;
  assign T1665 = T1671 ? readValueBankFifo : T1666;
  assign T1666 = T1667 ? readValueBankFifo : 32'h0;
  assign T1667 = T420 & T1668;
  assign T1668 = T1669[5'h13:5'h13];
  assign T1669 = 1'h1 << T1670;
  assign T1670 = T3133;
  assign T3133 = {2'h0, portId};
  assign T1671 = T423 & T1668;
  assign T1672 = T1681 | T1673;
  assign T1673 = bankToPort_3_19;
  assign bankToPort_3_19 = T1674;
  assign T1674 = T1680 ? readValueBankFifo : T1675;
  assign T1675 = T1676 ? readValueBankFifo : 32'h0;
  assign T1676 = T415 & T1677;
  assign T1677 = T1678[5'h13:5'h13];
  assign T1678 = 1'h1 << T1679;
  assign T1679 = T3134;
  assign T3134 = {2'h0, portId};
  assign T1680 = T418 & T1677;
  assign T1681 = T1690 | T1682;
  assign T1682 = bankToPort_2_19;
  assign bankToPort_2_19 = T1683;
  assign T1683 = T1689 ? readValueBankFifo : T1684;
  assign T1684 = T1685 ? readValueBankFifo : 32'h0;
  assign T1685 = T410 & T1686;
  assign T1686 = T1687[5'h13:5'h13];
  assign T1687 = 1'h1 << T1688;
  assign T1688 = T3135;
  assign T3135 = {2'h0, portId};
  assign T1689 = T413 & T1686;
  assign T1690 = T1699 | T1691;
  assign T1691 = bankToPort_1_19;
  assign bankToPort_1_19 = T1692;
  assign T1692 = T1698 ? readValueBankFifo : T1693;
  assign T1693 = T1694 ? readValueBankFifo : 32'h0;
  assign T1694 = T405 & T1695;
  assign T1695 = T1696[5'h13:5'h13];
  assign T1696 = 1'h1 << T1697;
  assign T1697 = T3136;
  assign T3136 = {2'h0, portId};
  assign T1698 = T408 & T1695;
  assign T1699 = 32'h1 | T1700;
  assign T1700 = bankToPort_0_19;
  assign bankToPort_0_19 = T1701;
  assign T1701 = T1707 ? readValueBankFifo : T1702;
  assign T1702 = T1703 ? readValueBankFifo : 32'h0;
  assign T1703 = T402 & T1704;
  assign T1704 = T1705[5'h13:5'h13];
  assign T1705 = 1'h1 << T1706;
  assign T1706 = T3137;
  assign T3137 = {2'h0, portId};
  assign T1707 = T500 & T1704;
  assign T1708 = T1509 ^ 1'h1;
  assign T1709 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1710 = T1711 ? 1'h1 : 1'h0;
  assign T1711 = T1453 & fifo_38_io_enqRdy;
  assign T1712 = seqLevelDoneReg2 ? fifo_18_io_enqRdy : 1'h0;
  assign T1713 = T1711 ? T1714 : T1714;
  assign T1714 = T1715;
  assign T1715 = T1773 ? 32'h0 : T1716;
  assign T1716 = T1453 ? T1717 : 32'h0;
  assign T1717 = T1724 | T1718;
  assign T1718 = bankToPort_7_18;
  assign bankToPort_7_18 = T1719;
  assign T1719 = T1723 ? readValueBankFifo : T1720;
  assign T1720 = T1721 ? readValueBankFifo : 32'h0;
  assign T1721 = T269 & T1722;
  assign T1722 = T1627[5'h12:5'h12];
  assign T1723 = T436 & T1722;
  assign T1724 = T1731 | T1725;
  assign T1725 = bankToPort_6_18;
  assign bankToPort_6_18 = T1726;
  assign T1726 = T1730 ? readValueBankFifo : T1727;
  assign T1727 = T1728 ? readValueBankFifo : 32'h0;
  assign T1728 = T430 & T1729;
  assign T1729 = T1651[5'h12:5'h12];
  assign T1730 = T433 & T1729;
  assign T1731 = T1738 | T1732;
  assign T1732 = bankToPort_5_18;
  assign bankToPort_5_18 = T1733;
  assign T1733 = T1737 ? readValueBankFifo : T1734;
  assign T1734 = T1735 ? readValueBankFifo : 32'h0;
  assign T1735 = T425 & T1736;
  assign T1736 = T1660[5'h12:5'h12];
  assign T1737 = T428 & T1736;
  assign T1738 = T1745 | T1739;
  assign T1739 = bankToPort_4_18;
  assign bankToPort_4_18 = T1740;
  assign T1740 = T1744 ? readValueBankFifo : T1741;
  assign T1741 = T1742 ? readValueBankFifo : 32'h0;
  assign T1742 = T420 & T1743;
  assign T1743 = T1669[5'h12:5'h12];
  assign T1744 = T423 & T1743;
  assign T1745 = T1752 | T1746;
  assign T1746 = bankToPort_3_18;
  assign bankToPort_3_18 = T1747;
  assign T1747 = T1751 ? readValueBankFifo : T1748;
  assign T1748 = T1749 ? readValueBankFifo : 32'h0;
  assign T1749 = T415 & T1750;
  assign T1750 = T1678[5'h12:5'h12];
  assign T1751 = T418 & T1750;
  assign T1752 = T1759 | T1753;
  assign T1753 = bankToPort_2_18;
  assign bankToPort_2_18 = T1754;
  assign T1754 = T1758 ? readValueBankFifo : T1755;
  assign T1755 = T1756 ? readValueBankFifo : 32'h0;
  assign T1756 = T410 & T1757;
  assign T1757 = T1687[5'h12:5'h12];
  assign T1758 = T413 & T1757;
  assign T1759 = T1766 | T1760;
  assign T1760 = bankToPort_1_18;
  assign bankToPort_1_18 = T1761;
  assign T1761 = T1765 ? readValueBankFifo : T1762;
  assign T1762 = T1763 ? readValueBankFifo : 32'h0;
  assign T1763 = T405 & T1764;
  assign T1764 = T1696[5'h12:5'h12];
  assign T1765 = T408 & T1764;
  assign T1766 = 32'h1 | T1767;
  assign T1767 = bankToPort_0_18;
  assign bankToPort_0_18 = T1768;
  assign T1768 = T1772 ? readValueBankFifo : T1769;
  assign T1769 = T1770 ? readValueBankFifo : 32'h0;
  assign T1770 = T402 & T1771;
  assign T1771 = T1705[5'h12:5'h12];
  assign T1772 = T500 & T1771;
  assign T1773 = T1453 ^ 1'h1;
  assign T1774 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1775 = T1776 ? 1'h1 : 1'h0;
  assign T1776 = T1397 & fifo_37_io_enqRdy;
  assign T1777 = seqLevelDoneReg2 ? fifo_17_io_enqRdy : 1'h0;
  assign T1778 = T1776 ? T1779 : T1779;
  assign T1779 = T1780;
  assign T1780 = T1838 ? 32'h0 : T1781;
  assign T1781 = T1397 ? T1782 : 32'h0;
  assign T1782 = T1789 | T1783;
  assign T1783 = bankToPort_7_17;
  assign bankToPort_7_17 = T1784;
  assign T1784 = T1788 ? readValueBankFifo : T1785;
  assign T1785 = T1786 ? readValueBankFifo : 32'h0;
  assign T1786 = T269 & T1787;
  assign T1787 = T1627[5'h11:5'h11];
  assign T1788 = T436 & T1787;
  assign T1789 = T1796 | T1790;
  assign T1790 = bankToPort_6_17;
  assign bankToPort_6_17 = T1791;
  assign T1791 = T1795 ? readValueBankFifo : T1792;
  assign T1792 = T1793 ? readValueBankFifo : 32'h0;
  assign T1793 = T430 & T1794;
  assign T1794 = T1651[5'h11:5'h11];
  assign T1795 = T433 & T1794;
  assign T1796 = T1803 | T1797;
  assign T1797 = bankToPort_5_17;
  assign bankToPort_5_17 = T1798;
  assign T1798 = T1802 ? readValueBankFifo : T1799;
  assign T1799 = T1800 ? readValueBankFifo : 32'h0;
  assign T1800 = T425 & T1801;
  assign T1801 = T1660[5'h11:5'h11];
  assign T1802 = T428 & T1801;
  assign T1803 = T1810 | T1804;
  assign T1804 = bankToPort_4_17;
  assign bankToPort_4_17 = T1805;
  assign T1805 = T1809 ? readValueBankFifo : T1806;
  assign T1806 = T1807 ? readValueBankFifo : 32'h0;
  assign T1807 = T420 & T1808;
  assign T1808 = T1669[5'h11:5'h11];
  assign T1809 = T423 & T1808;
  assign T1810 = T1817 | T1811;
  assign T1811 = bankToPort_3_17;
  assign bankToPort_3_17 = T1812;
  assign T1812 = T1816 ? readValueBankFifo : T1813;
  assign T1813 = T1814 ? readValueBankFifo : 32'h0;
  assign T1814 = T415 & T1815;
  assign T1815 = T1678[5'h11:5'h11];
  assign T1816 = T418 & T1815;
  assign T1817 = T1824 | T1818;
  assign T1818 = bankToPort_2_17;
  assign bankToPort_2_17 = T1819;
  assign T1819 = T1823 ? readValueBankFifo : T1820;
  assign T1820 = T1821 ? readValueBankFifo : 32'h0;
  assign T1821 = T410 & T1822;
  assign T1822 = T1687[5'h11:5'h11];
  assign T1823 = T413 & T1822;
  assign T1824 = T1831 | T1825;
  assign T1825 = bankToPort_1_17;
  assign bankToPort_1_17 = T1826;
  assign T1826 = T1830 ? readValueBankFifo : T1827;
  assign T1827 = T1828 ? readValueBankFifo : 32'h0;
  assign T1828 = T405 & T1829;
  assign T1829 = T1696[5'h11:5'h11];
  assign T1830 = T408 & T1829;
  assign T1831 = 32'h1 | T1832;
  assign T1832 = bankToPort_0_17;
  assign bankToPort_0_17 = T1833;
  assign T1833 = T1837 ? readValueBankFifo : T1834;
  assign T1834 = T1835 ? readValueBankFifo : 32'h0;
  assign T1835 = T402 & T1836;
  assign T1836 = T1705[5'h11:5'h11];
  assign T1837 = T500 & T1836;
  assign T1838 = T1397 ^ 1'h1;
  assign T1839 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1840 = T1841 ? 1'h1 : 1'h0;
  assign T1841 = T1341 & fifo_36_io_enqRdy;
  assign T1842 = seqLevelDoneReg2 ? fifo_16_io_enqRdy : 1'h0;
  assign T1843 = T1841 ? T1844 : T1844;
  assign T1844 = T1845;
  assign T1845 = T1903 ? 32'h0 : T1846;
  assign T1846 = T1341 ? T1847 : 32'h0;
  assign T1847 = T1854 | T1848;
  assign T1848 = bankToPort_7_16;
  assign bankToPort_7_16 = T1849;
  assign T1849 = T1853 ? readValueBankFifo : T1850;
  assign T1850 = T1851 ? readValueBankFifo : 32'h0;
  assign T1851 = T269 & T1852;
  assign T1852 = T1627[5'h10:5'h10];
  assign T1853 = T436 & T1852;
  assign T1854 = T1861 | T1855;
  assign T1855 = bankToPort_6_16;
  assign bankToPort_6_16 = T1856;
  assign T1856 = T1860 ? readValueBankFifo : T1857;
  assign T1857 = T1858 ? readValueBankFifo : 32'h0;
  assign T1858 = T430 & T1859;
  assign T1859 = T1651[5'h10:5'h10];
  assign T1860 = T433 & T1859;
  assign T1861 = T1868 | T1862;
  assign T1862 = bankToPort_5_16;
  assign bankToPort_5_16 = T1863;
  assign T1863 = T1867 ? readValueBankFifo : T1864;
  assign T1864 = T1865 ? readValueBankFifo : 32'h0;
  assign T1865 = T425 & T1866;
  assign T1866 = T1660[5'h10:5'h10];
  assign T1867 = T428 & T1866;
  assign T1868 = T1875 | T1869;
  assign T1869 = bankToPort_4_16;
  assign bankToPort_4_16 = T1870;
  assign T1870 = T1874 ? readValueBankFifo : T1871;
  assign T1871 = T1872 ? readValueBankFifo : 32'h0;
  assign T1872 = T420 & T1873;
  assign T1873 = T1669[5'h10:5'h10];
  assign T1874 = T423 & T1873;
  assign T1875 = T1882 | T1876;
  assign T1876 = bankToPort_3_16;
  assign bankToPort_3_16 = T1877;
  assign T1877 = T1881 ? readValueBankFifo : T1878;
  assign T1878 = T1879 ? readValueBankFifo : 32'h0;
  assign T1879 = T415 & T1880;
  assign T1880 = T1678[5'h10:5'h10];
  assign T1881 = T418 & T1880;
  assign T1882 = T1889 | T1883;
  assign T1883 = bankToPort_2_16;
  assign bankToPort_2_16 = T1884;
  assign T1884 = T1888 ? readValueBankFifo : T1885;
  assign T1885 = T1886 ? readValueBankFifo : 32'h0;
  assign T1886 = T410 & T1887;
  assign T1887 = T1687[5'h10:5'h10];
  assign T1888 = T413 & T1887;
  assign T1889 = T1896 | T1890;
  assign T1890 = bankToPort_1_16;
  assign bankToPort_1_16 = T1891;
  assign T1891 = T1895 ? readValueBankFifo : T1892;
  assign T1892 = T1893 ? readValueBankFifo : 32'h0;
  assign T1893 = T405 & T1894;
  assign T1894 = T1696[5'h10:5'h10];
  assign T1895 = T408 & T1894;
  assign T1896 = 32'h1 | T1897;
  assign T1897 = bankToPort_0_16;
  assign bankToPort_0_16 = T1898;
  assign T1898 = T1902 ? readValueBankFifo : T1899;
  assign T1899 = T1900 ? readValueBankFifo : 32'h0;
  assign T1900 = T402 & T1901;
  assign T1901 = T1705[5'h10:5'h10];
  assign T1902 = T500 & T1901;
  assign T1903 = T1341 ^ 1'h1;
  assign T1904 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1905 = T1906 ? 1'h1 : 1'h0;
  assign T1906 = T1285 & fifo_35_io_enqRdy;
  assign T1907 = seqLevelDoneReg2 ? fifo_15_io_enqRdy : 1'h0;
  assign T1908 = T1906 ? T1909 : T1909;
  assign T1909 = T1910;
  assign T1910 = T1968 ? 32'h0 : T1911;
  assign T1911 = T1285 ? T1912 : 32'h0;
  assign T1912 = T1919 | T1913;
  assign T1913 = bankToPort_7_15;
  assign bankToPort_7_15 = T1914;
  assign T1914 = T1918 ? readValueBankFifo : T1915;
  assign T1915 = T1916 ? readValueBankFifo : 32'h0;
  assign T1916 = T269 & T1917;
  assign T1917 = T1627[4'hf:4'hf];
  assign T1918 = T436 & T1917;
  assign T1919 = T1926 | T1920;
  assign T1920 = bankToPort_6_15;
  assign bankToPort_6_15 = T1921;
  assign T1921 = T1925 ? readValueBankFifo : T1922;
  assign T1922 = T1923 ? readValueBankFifo : 32'h0;
  assign T1923 = T430 & T1924;
  assign T1924 = T1651[4'hf:4'hf];
  assign T1925 = T433 & T1924;
  assign T1926 = T1933 | T1927;
  assign T1927 = bankToPort_5_15;
  assign bankToPort_5_15 = T1928;
  assign T1928 = T1932 ? readValueBankFifo : T1929;
  assign T1929 = T1930 ? readValueBankFifo : 32'h0;
  assign T1930 = T425 & T1931;
  assign T1931 = T1660[4'hf:4'hf];
  assign T1932 = T428 & T1931;
  assign T1933 = T1940 | T1934;
  assign T1934 = bankToPort_4_15;
  assign bankToPort_4_15 = T1935;
  assign T1935 = T1939 ? readValueBankFifo : T1936;
  assign T1936 = T1937 ? readValueBankFifo : 32'h0;
  assign T1937 = T420 & T1938;
  assign T1938 = T1669[4'hf:4'hf];
  assign T1939 = T423 & T1938;
  assign T1940 = T1947 | T1941;
  assign T1941 = bankToPort_3_15;
  assign bankToPort_3_15 = T1942;
  assign T1942 = T1946 ? readValueBankFifo : T1943;
  assign T1943 = T1944 ? readValueBankFifo : 32'h0;
  assign T1944 = T415 & T1945;
  assign T1945 = T1678[4'hf:4'hf];
  assign T1946 = T418 & T1945;
  assign T1947 = T1954 | T1948;
  assign T1948 = bankToPort_2_15;
  assign bankToPort_2_15 = T1949;
  assign T1949 = T1953 ? readValueBankFifo : T1950;
  assign T1950 = T1951 ? readValueBankFifo : 32'h0;
  assign T1951 = T410 & T1952;
  assign T1952 = T1687[4'hf:4'hf];
  assign T1953 = T413 & T1952;
  assign T1954 = T1961 | T1955;
  assign T1955 = bankToPort_1_15;
  assign bankToPort_1_15 = T1956;
  assign T1956 = T1960 ? readValueBankFifo : T1957;
  assign T1957 = T1958 ? readValueBankFifo : 32'h0;
  assign T1958 = T405 & T1959;
  assign T1959 = T1696[4'hf:4'hf];
  assign T1960 = T408 & T1959;
  assign T1961 = 32'h1 | T1962;
  assign T1962 = bankToPort_0_15;
  assign bankToPort_0_15 = T1963;
  assign T1963 = T1967 ? readValueBankFifo : T1964;
  assign T1964 = T1965 ? readValueBankFifo : 32'h0;
  assign T1965 = T402 & T1966;
  assign T1966 = T1705[4'hf:4'hf];
  assign T1967 = T500 & T1966;
  assign T1968 = T1285 ^ 1'h1;
  assign T1969 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1970 = T1971 ? 1'h1 : 1'h0;
  assign T1971 = T1229 & fifo_34_io_enqRdy;
  assign T1972 = seqLevelDoneReg2 ? fifo_14_io_enqRdy : 1'h0;
  assign T1973 = T1971 ? T1974 : T1974;
  assign T1974 = T1975;
  assign T1975 = T2033 ? 32'h0 : T1976;
  assign T1976 = T1229 ? T1977 : 32'h0;
  assign T1977 = T1984 | T1978;
  assign T1978 = bankToPort_7_14;
  assign bankToPort_7_14 = T1979;
  assign T1979 = T1983 ? readValueBankFifo : T1980;
  assign T1980 = T1981 ? readValueBankFifo : 32'h0;
  assign T1981 = T269 & T1982;
  assign T1982 = T1627[4'he:4'he];
  assign T1983 = T436 & T1982;
  assign T1984 = T1991 | T1985;
  assign T1985 = bankToPort_6_14;
  assign bankToPort_6_14 = T1986;
  assign T1986 = T1990 ? readValueBankFifo : T1987;
  assign T1987 = T1988 ? readValueBankFifo : 32'h0;
  assign T1988 = T430 & T1989;
  assign T1989 = T1651[4'he:4'he];
  assign T1990 = T433 & T1989;
  assign T1991 = T1998 | T1992;
  assign T1992 = bankToPort_5_14;
  assign bankToPort_5_14 = T1993;
  assign T1993 = T1997 ? readValueBankFifo : T1994;
  assign T1994 = T1995 ? readValueBankFifo : 32'h0;
  assign T1995 = T425 & T1996;
  assign T1996 = T1660[4'he:4'he];
  assign T1997 = T428 & T1996;
  assign T1998 = T2005 | T1999;
  assign T1999 = bankToPort_4_14;
  assign bankToPort_4_14 = T2000;
  assign T2000 = T2004 ? readValueBankFifo : T2001;
  assign T2001 = T2002 ? readValueBankFifo : 32'h0;
  assign T2002 = T420 & T2003;
  assign T2003 = T1669[4'he:4'he];
  assign T2004 = T423 & T2003;
  assign T2005 = T2012 | T2006;
  assign T2006 = bankToPort_3_14;
  assign bankToPort_3_14 = T2007;
  assign T2007 = T2011 ? readValueBankFifo : T2008;
  assign T2008 = T2009 ? readValueBankFifo : 32'h0;
  assign T2009 = T415 & T2010;
  assign T2010 = T1678[4'he:4'he];
  assign T2011 = T418 & T2010;
  assign T2012 = T2019 | T2013;
  assign T2013 = bankToPort_2_14;
  assign bankToPort_2_14 = T2014;
  assign T2014 = T2018 ? readValueBankFifo : T2015;
  assign T2015 = T2016 ? readValueBankFifo : 32'h0;
  assign T2016 = T410 & T2017;
  assign T2017 = T1687[4'he:4'he];
  assign T2018 = T413 & T2017;
  assign T2019 = T2026 | T2020;
  assign T2020 = bankToPort_1_14;
  assign bankToPort_1_14 = T2021;
  assign T2021 = T2025 ? readValueBankFifo : T2022;
  assign T2022 = T2023 ? readValueBankFifo : 32'h0;
  assign T2023 = T405 & T2024;
  assign T2024 = T1696[4'he:4'he];
  assign T2025 = T408 & T2024;
  assign T2026 = 32'h1 | T2027;
  assign T2027 = bankToPort_0_14;
  assign bankToPort_0_14 = T2028;
  assign T2028 = T2032 ? readValueBankFifo : T2029;
  assign T2029 = T2030 ? readValueBankFifo : 32'h0;
  assign T2030 = T402 & T2031;
  assign T2031 = T1705[4'he:4'he];
  assign T2032 = T500 & T2031;
  assign T2033 = T1229 ^ 1'h1;
  assign T2034 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2035 = T2036 ? 1'h1 : 1'h0;
  assign T2036 = T1173 & fifo_33_io_enqRdy;
  assign T2037 = seqLevelDoneReg2 ? fifo_13_io_enqRdy : 1'h0;
  assign T2038 = T2036 ? T2039 : T2039;
  assign T2039 = T2040;
  assign T2040 = T2098 ? 32'h0 : T2041;
  assign T2041 = T1173 ? T2042 : 32'h0;
  assign T2042 = T2049 | T2043;
  assign T2043 = bankToPort_7_13;
  assign bankToPort_7_13 = T2044;
  assign T2044 = T2048 ? readValueBankFifo : T2045;
  assign T2045 = T2046 ? readValueBankFifo : 32'h0;
  assign T2046 = T269 & T2047;
  assign T2047 = T1627[4'hd:4'hd];
  assign T2048 = T436 & T2047;
  assign T2049 = T2056 | T2050;
  assign T2050 = bankToPort_6_13;
  assign bankToPort_6_13 = T2051;
  assign T2051 = T2055 ? readValueBankFifo : T2052;
  assign T2052 = T2053 ? readValueBankFifo : 32'h0;
  assign T2053 = T430 & T2054;
  assign T2054 = T1651[4'hd:4'hd];
  assign T2055 = T433 & T2054;
  assign T2056 = T2063 | T2057;
  assign T2057 = bankToPort_5_13;
  assign bankToPort_5_13 = T2058;
  assign T2058 = T2062 ? readValueBankFifo : T2059;
  assign T2059 = T2060 ? readValueBankFifo : 32'h0;
  assign T2060 = T425 & T2061;
  assign T2061 = T1660[4'hd:4'hd];
  assign T2062 = T428 & T2061;
  assign T2063 = T2070 | T2064;
  assign T2064 = bankToPort_4_13;
  assign bankToPort_4_13 = T2065;
  assign T2065 = T2069 ? readValueBankFifo : T2066;
  assign T2066 = T2067 ? readValueBankFifo : 32'h0;
  assign T2067 = T420 & T2068;
  assign T2068 = T1669[4'hd:4'hd];
  assign T2069 = T423 & T2068;
  assign T2070 = T2077 | T2071;
  assign T2071 = bankToPort_3_13;
  assign bankToPort_3_13 = T2072;
  assign T2072 = T2076 ? readValueBankFifo : T2073;
  assign T2073 = T2074 ? readValueBankFifo : 32'h0;
  assign T2074 = T415 & T2075;
  assign T2075 = T1678[4'hd:4'hd];
  assign T2076 = T418 & T2075;
  assign T2077 = T2084 | T2078;
  assign T2078 = bankToPort_2_13;
  assign bankToPort_2_13 = T2079;
  assign T2079 = T2083 ? readValueBankFifo : T2080;
  assign T2080 = T2081 ? readValueBankFifo : 32'h0;
  assign T2081 = T410 & T2082;
  assign T2082 = T1687[4'hd:4'hd];
  assign T2083 = T413 & T2082;
  assign T2084 = T2091 | T2085;
  assign T2085 = bankToPort_1_13;
  assign bankToPort_1_13 = T2086;
  assign T2086 = T2090 ? readValueBankFifo : T2087;
  assign T2087 = T2088 ? readValueBankFifo : 32'h0;
  assign T2088 = T405 & T2089;
  assign T2089 = T1696[4'hd:4'hd];
  assign T2090 = T408 & T2089;
  assign T2091 = 32'h1 | T2092;
  assign T2092 = bankToPort_0_13;
  assign bankToPort_0_13 = T2093;
  assign T2093 = T2097 ? readValueBankFifo : T2094;
  assign T2094 = T2095 ? readValueBankFifo : 32'h0;
  assign T2095 = T402 & T2096;
  assign T2096 = T1705[4'hd:4'hd];
  assign T2097 = T500 & T2096;
  assign T2098 = T1173 ^ 1'h1;
  assign T2099 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2100 = T2101 ? 1'h1 : 1'h0;
  assign T2101 = T1117 & fifo_32_io_enqRdy;
  assign T2102 = seqLevelDoneReg2 ? fifo_12_io_enqRdy : 1'h0;
  assign T2103 = T2101 ? T2104 : T2104;
  assign T2104 = T2105;
  assign T2105 = T2163 ? 32'h0 : T2106;
  assign T2106 = T1117 ? T2107 : 32'h0;
  assign T2107 = T2114 | T2108;
  assign T2108 = bankToPort_7_12;
  assign bankToPort_7_12 = T2109;
  assign T2109 = T2113 ? readValueBankFifo : T2110;
  assign T2110 = T2111 ? readValueBankFifo : 32'h0;
  assign T2111 = T269 & T2112;
  assign T2112 = T1627[4'hc:4'hc];
  assign T2113 = T436 & T2112;
  assign T2114 = T2121 | T2115;
  assign T2115 = bankToPort_6_12;
  assign bankToPort_6_12 = T2116;
  assign T2116 = T2120 ? readValueBankFifo : T2117;
  assign T2117 = T2118 ? readValueBankFifo : 32'h0;
  assign T2118 = T430 & T2119;
  assign T2119 = T1651[4'hc:4'hc];
  assign T2120 = T433 & T2119;
  assign T2121 = T2128 | T2122;
  assign T2122 = bankToPort_5_12;
  assign bankToPort_5_12 = T2123;
  assign T2123 = T2127 ? readValueBankFifo : T2124;
  assign T2124 = T2125 ? readValueBankFifo : 32'h0;
  assign T2125 = T425 & T2126;
  assign T2126 = T1660[4'hc:4'hc];
  assign T2127 = T428 & T2126;
  assign T2128 = T2135 | T2129;
  assign T2129 = bankToPort_4_12;
  assign bankToPort_4_12 = T2130;
  assign T2130 = T2134 ? readValueBankFifo : T2131;
  assign T2131 = T2132 ? readValueBankFifo : 32'h0;
  assign T2132 = T420 & T2133;
  assign T2133 = T1669[4'hc:4'hc];
  assign T2134 = T423 & T2133;
  assign T2135 = T2142 | T2136;
  assign T2136 = bankToPort_3_12;
  assign bankToPort_3_12 = T2137;
  assign T2137 = T2141 ? readValueBankFifo : T2138;
  assign T2138 = T2139 ? readValueBankFifo : 32'h0;
  assign T2139 = T415 & T2140;
  assign T2140 = T1678[4'hc:4'hc];
  assign T2141 = T418 & T2140;
  assign T2142 = T2149 | T2143;
  assign T2143 = bankToPort_2_12;
  assign bankToPort_2_12 = T2144;
  assign T2144 = T2148 ? readValueBankFifo : T2145;
  assign T2145 = T2146 ? readValueBankFifo : 32'h0;
  assign T2146 = T410 & T2147;
  assign T2147 = T1687[4'hc:4'hc];
  assign T2148 = T413 & T2147;
  assign T2149 = T2156 | T2150;
  assign T2150 = bankToPort_1_12;
  assign bankToPort_1_12 = T2151;
  assign T2151 = T2155 ? readValueBankFifo : T2152;
  assign T2152 = T2153 ? readValueBankFifo : 32'h0;
  assign T2153 = T405 & T2154;
  assign T2154 = T1696[4'hc:4'hc];
  assign T2155 = T408 & T2154;
  assign T2156 = 32'h1 | T2157;
  assign T2157 = bankToPort_0_12;
  assign bankToPort_0_12 = T2158;
  assign T2158 = T2162 ? readValueBankFifo : T2159;
  assign T2159 = T2160 ? readValueBankFifo : 32'h0;
  assign T2160 = T402 & T2161;
  assign T2161 = T1705[4'hc:4'hc];
  assign T2162 = T500 & T2161;
  assign T2163 = T1117 ^ 1'h1;
  assign T2164 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2165 = T2166 ? 1'h1 : 1'h0;
  assign T2166 = T1061 & fifo_31_io_enqRdy;
  assign T2167 = seqLevelDoneReg2 ? fifo_11_io_enqRdy : 1'h0;
  assign T2168 = T2166 ? T2169 : T2169;
  assign T2169 = T2170;
  assign T2170 = T2228 ? 32'h0 : T2171;
  assign T2171 = T1061 ? T2172 : 32'h0;
  assign T2172 = T2179 | T2173;
  assign T2173 = bankToPort_7_11;
  assign bankToPort_7_11 = T2174;
  assign T2174 = T2178 ? readValueBankFifo : T2175;
  assign T2175 = T2176 ? readValueBankFifo : 32'h0;
  assign T2176 = T269 & T2177;
  assign T2177 = T1627[4'hb:4'hb];
  assign T2178 = T436 & T2177;
  assign T2179 = T2186 | T2180;
  assign T2180 = bankToPort_6_11;
  assign bankToPort_6_11 = T2181;
  assign T2181 = T2185 ? readValueBankFifo : T2182;
  assign T2182 = T2183 ? readValueBankFifo : 32'h0;
  assign T2183 = T430 & T2184;
  assign T2184 = T1651[4'hb:4'hb];
  assign T2185 = T433 & T2184;
  assign T2186 = T2193 | T2187;
  assign T2187 = bankToPort_5_11;
  assign bankToPort_5_11 = T2188;
  assign T2188 = T2192 ? readValueBankFifo : T2189;
  assign T2189 = T2190 ? readValueBankFifo : 32'h0;
  assign T2190 = T425 & T2191;
  assign T2191 = T1660[4'hb:4'hb];
  assign T2192 = T428 & T2191;
  assign T2193 = T2200 | T2194;
  assign T2194 = bankToPort_4_11;
  assign bankToPort_4_11 = T2195;
  assign T2195 = T2199 ? readValueBankFifo : T2196;
  assign T2196 = T2197 ? readValueBankFifo : 32'h0;
  assign T2197 = T420 & T2198;
  assign T2198 = T1669[4'hb:4'hb];
  assign T2199 = T423 & T2198;
  assign T2200 = T2207 | T2201;
  assign T2201 = bankToPort_3_11;
  assign bankToPort_3_11 = T2202;
  assign T2202 = T2206 ? readValueBankFifo : T2203;
  assign T2203 = T2204 ? readValueBankFifo : 32'h0;
  assign T2204 = T415 & T2205;
  assign T2205 = T1678[4'hb:4'hb];
  assign T2206 = T418 & T2205;
  assign T2207 = T2214 | T2208;
  assign T2208 = bankToPort_2_11;
  assign bankToPort_2_11 = T2209;
  assign T2209 = T2213 ? readValueBankFifo : T2210;
  assign T2210 = T2211 ? readValueBankFifo : 32'h0;
  assign T2211 = T410 & T2212;
  assign T2212 = T1687[4'hb:4'hb];
  assign T2213 = T413 & T2212;
  assign T2214 = T2221 | T2215;
  assign T2215 = bankToPort_1_11;
  assign bankToPort_1_11 = T2216;
  assign T2216 = T2220 ? readValueBankFifo : T2217;
  assign T2217 = T2218 ? readValueBankFifo : 32'h0;
  assign T2218 = T405 & T2219;
  assign T2219 = T1696[4'hb:4'hb];
  assign T2220 = T408 & T2219;
  assign T2221 = 32'h1 | T2222;
  assign T2222 = bankToPort_0_11;
  assign bankToPort_0_11 = T2223;
  assign T2223 = T2227 ? readValueBankFifo : T2224;
  assign T2224 = T2225 ? readValueBankFifo : 32'h0;
  assign T2225 = T402 & T2226;
  assign T2226 = T1705[4'hb:4'hb];
  assign T2227 = T500 & T2226;
  assign T2228 = T1061 ^ 1'h1;
  assign T2229 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2230 = T2231 ? 1'h1 : 1'h0;
  assign T2231 = T1005 & fifo_30_io_enqRdy;
  assign T2232 = seqLevelDoneReg2 ? fifo_10_io_enqRdy : 1'h0;
  assign T2233 = T2231 ? T2234 : T2234;
  assign T2234 = T2235;
  assign T2235 = T2293 ? 32'h0 : T2236;
  assign T2236 = T1005 ? T2237 : 32'h0;
  assign T2237 = T2244 | T2238;
  assign T2238 = bankToPort_7_10;
  assign bankToPort_7_10 = T2239;
  assign T2239 = T2243 ? readValueBankFifo : T2240;
  assign T2240 = T2241 ? readValueBankFifo : 32'h0;
  assign T2241 = T269 & T2242;
  assign T2242 = T1627[4'ha:4'ha];
  assign T2243 = T436 & T2242;
  assign T2244 = T2251 | T2245;
  assign T2245 = bankToPort_6_10;
  assign bankToPort_6_10 = T2246;
  assign T2246 = T2250 ? readValueBankFifo : T2247;
  assign T2247 = T2248 ? readValueBankFifo : 32'h0;
  assign T2248 = T430 & T2249;
  assign T2249 = T1651[4'ha:4'ha];
  assign T2250 = T433 & T2249;
  assign T2251 = T2258 | T2252;
  assign T2252 = bankToPort_5_10;
  assign bankToPort_5_10 = T2253;
  assign T2253 = T2257 ? readValueBankFifo : T2254;
  assign T2254 = T2255 ? readValueBankFifo : 32'h0;
  assign T2255 = T425 & T2256;
  assign T2256 = T1660[4'ha:4'ha];
  assign T2257 = T428 & T2256;
  assign T2258 = T2265 | T2259;
  assign T2259 = bankToPort_4_10;
  assign bankToPort_4_10 = T2260;
  assign T2260 = T2264 ? readValueBankFifo : T2261;
  assign T2261 = T2262 ? readValueBankFifo : 32'h0;
  assign T2262 = T420 & T2263;
  assign T2263 = T1669[4'ha:4'ha];
  assign T2264 = T423 & T2263;
  assign T2265 = T2272 | T2266;
  assign T2266 = bankToPort_3_10;
  assign bankToPort_3_10 = T2267;
  assign T2267 = T2271 ? readValueBankFifo : T2268;
  assign T2268 = T2269 ? readValueBankFifo : 32'h0;
  assign T2269 = T415 & T2270;
  assign T2270 = T1678[4'ha:4'ha];
  assign T2271 = T418 & T2270;
  assign T2272 = T2279 | T2273;
  assign T2273 = bankToPort_2_10;
  assign bankToPort_2_10 = T2274;
  assign T2274 = T2278 ? readValueBankFifo : T2275;
  assign T2275 = T2276 ? readValueBankFifo : 32'h0;
  assign T2276 = T410 & T2277;
  assign T2277 = T1687[4'ha:4'ha];
  assign T2278 = T413 & T2277;
  assign T2279 = T2286 | T2280;
  assign T2280 = bankToPort_1_10;
  assign bankToPort_1_10 = T2281;
  assign T2281 = T2285 ? readValueBankFifo : T2282;
  assign T2282 = T2283 ? readValueBankFifo : 32'h0;
  assign T2283 = T405 & T2284;
  assign T2284 = T1696[4'ha:4'ha];
  assign T2285 = T408 & T2284;
  assign T2286 = 32'h1 | T2287;
  assign T2287 = bankToPort_0_10;
  assign bankToPort_0_10 = T2288;
  assign T2288 = T2292 ? readValueBankFifo : T2289;
  assign T2289 = T2290 ? readValueBankFifo : 32'h0;
  assign T2290 = T402 & T2291;
  assign T2291 = T1705[4'ha:4'ha];
  assign T2292 = T500 & T2291;
  assign T2293 = T1005 ^ 1'h1;
  assign T2294 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2295 = T2296 ? 1'h1 : 1'h0;
  assign T2296 = T949 & fifo_29_io_enqRdy;
  assign T2297 = seqLevelDoneReg2 ? fifo_9_io_enqRdy : 1'h0;
  assign T2298 = T2296 ? T2299 : T2299;
  assign T2299 = T2300;
  assign T2300 = T2358 ? 32'h0 : T2301;
  assign T2301 = T949 ? T2302 : 32'h0;
  assign T2302 = T2309 | T2303;
  assign T2303 = bankToPort_7_9;
  assign bankToPort_7_9 = T2304;
  assign T2304 = T2308 ? readValueBankFifo : T2305;
  assign T2305 = T2306 ? readValueBankFifo : 32'h0;
  assign T2306 = T269 & T2307;
  assign T2307 = T1627[4'h9:4'h9];
  assign T2308 = T436 & T2307;
  assign T2309 = T2316 | T2310;
  assign T2310 = bankToPort_6_9;
  assign bankToPort_6_9 = T2311;
  assign T2311 = T2315 ? readValueBankFifo : T2312;
  assign T2312 = T2313 ? readValueBankFifo : 32'h0;
  assign T2313 = T430 & T2314;
  assign T2314 = T1651[4'h9:4'h9];
  assign T2315 = T433 & T2314;
  assign T2316 = T2323 | T2317;
  assign T2317 = bankToPort_5_9;
  assign bankToPort_5_9 = T2318;
  assign T2318 = T2322 ? readValueBankFifo : T2319;
  assign T2319 = T2320 ? readValueBankFifo : 32'h0;
  assign T2320 = T425 & T2321;
  assign T2321 = T1660[4'h9:4'h9];
  assign T2322 = T428 & T2321;
  assign T2323 = T2330 | T2324;
  assign T2324 = bankToPort_4_9;
  assign bankToPort_4_9 = T2325;
  assign T2325 = T2329 ? readValueBankFifo : T2326;
  assign T2326 = T2327 ? readValueBankFifo : 32'h0;
  assign T2327 = T420 & T2328;
  assign T2328 = T1669[4'h9:4'h9];
  assign T2329 = T423 & T2328;
  assign T2330 = T2337 | T2331;
  assign T2331 = bankToPort_3_9;
  assign bankToPort_3_9 = T2332;
  assign T2332 = T2336 ? readValueBankFifo : T2333;
  assign T2333 = T2334 ? readValueBankFifo : 32'h0;
  assign T2334 = T415 & T2335;
  assign T2335 = T1678[4'h9:4'h9];
  assign T2336 = T418 & T2335;
  assign T2337 = T2344 | T2338;
  assign T2338 = bankToPort_2_9;
  assign bankToPort_2_9 = T2339;
  assign T2339 = T2343 ? readValueBankFifo : T2340;
  assign T2340 = T2341 ? readValueBankFifo : 32'h0;
  assign T2341 = T410 & T2342;
  assign T2342 = T1687[4'h9:4'h9];
  assign T2343 = T413 & T2342;
  assign T2344 = T2351 | T2345;
  assign T2345 = bankToPort_1_9;
  assign bankToPort_1_9 = T2346;
  assign T2346 = T2350 ? readValueBankFifo : T2347;
  assign T2347 = T2348 ? readValueBankFifo : 32'h0;
  assign T2348 = T405 & T2349;
  assign T2349 = T1696[4'h9:4'h9];
  assign T2350 = T408 & T2349;
  assign T2351 = 32'h1 | T2352;
  assign T2352 = bankToPort_0_9;
  assign bankToPort_0_9 = T2353;
  assign T2353 = T2357 ? readValueBankFifo : T2354;
  assign T2354 = T2355 ? readValueBankFifo : 32'h0;
  assign T2355 = T402 & T2356;
  assign T2356 = T1705[4'h9:4'h9];
  assign T2357 = T500 & T2356;
  assign T2358 = T949 ^ 1'h1;
  assign T2359 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2360 = T2361 ? 1'h1 : 1'h0;
  assign T2361 = T893 & fifo_28_io_enqRdy;
  assign T2362 = seqLevelDoneReg2 ? fifo_8_io_enqRdy : 1'h0;
  assign T2363 = T2361 ? T2364 : T2364;
  assign T2364 = T2365;
  assign T2365 = T2423 ? 32'h0 : T2366;
  assign T2366 = T893 ? T2367 : 32'h0;
  assign T2367 = T2374 | T2368;
  assign T2368 = bankToPort_7_8;
  assign bankToPort_7_8 = T2369;
  assign T2369 = T2373 ? readValueBankFifo : T2370;
  assign T2370 = T2371 ? readValueBankFifo : 32'h0;
  assign T2371 = T269 & T2372;
  assign T2372 = T1627[4'h8:4'h8];
  assign T2373 = T436 & T2372;
  assign T2374 = T2381 | T2375;
  assign T2375 = bankToPort_6_8;
  assign bankToPort_6_8 = T2376;
  assign T2376 = T2380 ? readValueBankFifo : T2377;
  assign T2377 = T2378 ? readValueBankFifo : 32'h0;
  assign T2378 = T430 & T2379;
  assign T2379 = T1651[4'h8:4'h8];
  assign T2380 = T433 & T2379;
  assign T2381 = T2388 | T2382;
  assign T2382 = bankToPort_5_8;
  assign bankToPort_5_8 = T2383;
  assign T2383 = T2387 ? readValueBankFifo : T2384;
  assign T2384 = T2385 ? readValueBankFifo : 32'h0;
  assign T2385 = T425 & T2386;
  assign T2386 = T1660[4'h8:4'h8];
  assign T2387 = T428 & T2386;
  assign T2388 = T2395 | T2389;
  assign T2389 = bankToPort_4_8;
  assign bankToPort_4_8 = T2390;
  assign T2390 = T2394 ? readValueBankFifo : T2391;
  assign T2391 = T2392 ? readValueBankFifo : 32'h0;
  assign T2392 = T420 & T2393;
  assign T2393 = T1669[4'h8:4'h8];
  assign T2394 = T423 & T2393;
  assign T2395 = T2402 | T2396;
  assign T2396 = bankToPort_3_8;
  assign bankToPort_3_8 = T2397;
  assign T2397 = T2401 ? readValueBankFifo : T2398;
  assign T2398 = T2399 ? readValueBankFifo : 32'h0;
  assign T2399 = T415 & T2400;
  assign T2400 = T1678[4'h8:4'h8];
  assign T2401 = T418 & T2400;
  assign T2402 = T2409 | T2403;
  assign T2403 = bankToPort_2_8;
  assign bankToPort_2_8 = T2404;
  assign T2404 = T2408 ? readValueBankFifo : T2405;
  assign T2405 = T2406 ? readValueBankFifo : 32'h0;
  assign T2406 = T410 & T2407;
  assign T2407 = T1687[4'h8:4'h8];
  assign T2408 = T413 & T2407;
  assign T2409 = T2416 | T2410;
  assign T2410 = bankToPort_1_8;
  assign bankToPort_1_8 = T2411;
  assign T2411 = T2415 ? readValueBankFifo : T2412;
  assign T2412 = T2413 ? readValueBankFifo : 32'h0;
  assign T2413 = T405 & T2414;
  assign T2414 = T1696[4'h8:4'h8];
  assign T2415 = T408 & T2414;
  assign T2416 = 32'h1 | T2417;
  assign T2417 = bankToPort_0_8;
  assign bankToPort_0_8 = T2418;
  assign T2418 = T2422 ? readValueBankFifo : T2419;
  assign T2419 = T2420 ? readValueBankFifo : 32'h0;
  assign T2420 = T402 & T2421;
  assign T2421 = T1705[4'h8:4'h8];
  assign T2422 = T500 & T2421;
  assign T2423 = T893 ^ 1'h1;
  assign T2424 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2425 = T2426 ? 1'h1 : 1'h0;
  assign T2426 = T837 & fifo_27_io_enqRdy;
  assign T2427 = seqLevelDoneReg2 ? fifo_7_io_enqRdy : 1'h0;
  assign T2428 = T2426 ? T2429 : T2429;
  assign T2429 = T2430;
  assign T2430 = T2488 ? 32'h0 : T2431;
  assign T2431 = T837 ? T2432 : 32'h0;
  assign T2432 = T2439 | T2433;
  assign T2433 = bankToPort_7_7;
  assign bankToPort_7_7 = T2434;
  assign T2434 = T2438 ? readValueBankFifo : T2435;
  assign T2435 = T2436 ? readValueBankFifo : 32'h0;
  assign T2436 = T269 & T2437;
  assign T2437 = T1627[3'h7:3'h7];
  assign T2438 = T436 & T2437;
  assign T2439 = T2446 | T2440;
  assign T2440 = bankToPort_6_7;
  assign bankToPort_6_7 = T2441;
  assign T2441 = T2445 ? readValueBankFifo : T2442;
  assign T2442 = T2443 ? readValueBankFifo : 32'h0;
  assign T2443 = T430 & T2444;
  assign T2444 = T1651[3'h7:3'h7];
  assign T2445 = T433 & T2444;
  assign T2446 = T2453 | T2447;
  assign T2447 = bankToPort_5_7;
  assign bankToPort_5_7 = T2448;
  assign T2448 = T2452 ? readValueBankFifo : T2449;
  assign T2449 = T2450 ? readValueBankFifo : 32'h0;
  assign T2450 = T425 & T2451;
  assign T2451 = T1660[3'h7:3'h7];
  assign T2452 = T428 & T2451;
  assign T2453 = T2460 | T2454;
  assign T2454 = bankToPort_4_7;
  assign bankToPort_4_7 = T2455;
  assign T2455 = T2459 ? readValueBankFifo : T2456;
  assign T2456 = T2457 ? readValueBankFifo : 32'h0;
  assign T2457 = T420 & T2458;
  assign T2458 = T1669[3'h7:3'h7];
  assign T2459 = T423 & T2458;
  assign T2460 = T2467 | T2461;
  assign T2461 = bankToPort_3_7;
  assign bankToPort_3_7 = T2462;
  assign T2462 = T2466 ? readValueBankFifo : T2463;
  assign T2463 = T2464 ? readValueBankFifo : 32'h0;
  assign T2464 = T415 & T2465;
  assign T2465 = T1678[3'h7:3'h7];
  assign T2466 = T418 & T2465;
  assign T2467 = T2474 | T2468;
  assign T2468 = bankToPort_2_7;
  assign bankToPort_2_7 = T2469;
  assign T2469 = T2473 ? readValueBankFifo : T2470;
  assign T2470 = T2471 ? readValueBankFifo : 32'h0;
  assign T2471 = T410 & T2472;
  assign T2472 = T1687[3'h7:3'h7];
  assign T2473 = T413 & T2472;
  assign T2474 = T2481 | T2475;
  assign T2475 = bankToPort_1_7;
  assign bankToPort_1_7 = T2476;
  assign T2476 = T2480 ? readValueBankFifo : T2477;
  assign T2477 = T2478 ? readValueBankFifo : 32'h0;
  assign T2478 = T405 & T2479;
  assign T2479 = T1696[3'h7:3'h7];
  assign T2480 = T408 & T2479;
  assign T2481 = 32'h1 | T2482;
  assign T2482 = bankToPort_0_7;
  assign bankToPort_0_7 = T2483;
  assign T2483 = T2487 ? readValueBankFifo : T2484;
  assign T2484 = T2485 ? readValueBankFifo : 32'h0;
  assign T2485 = T402 & T2486;
  assign T2486 = T1705[3'h7:3'h7];
  assign T2487 = T500 & T2486;
  assign T2488 = T837 ^ 1'h1;
  assign T2489 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2490 = T2491 ? 1'h1 : 1'h0;
  assign T2491 = T781 & fifo_26_io_enqRdy;
  assign T2492 = seqLevelDoneReg2 ? fifo_6_io_enqRdy : 1'h0;
  assign T2493 = T2491 ? T2494 : T2494;
  assign T2494 = T2495;
  assign T2495 = T2553 ? 32'h0 : T2496;
  assign T2496 = T781 ? T2497 : 32'h0;
  assign T2497 = T2504 | T2498;
  assign T2498 = bankToPort_7_6;
  assign bankToPort_7_6 = T2499;
  assign T2499 = T2503 ? readValueBankFifo : T2500;
  assign T2500 = T2501 ? readValueBankFifo : 32'h0;
  assign T2501 = T269 & T2502;
  assign T2502 = T1627[3'h6:3'h6];
  assign T2503 = T436 & T2502;
  assign T2504 = T2511 | T2505;
  assign T2505 = bankToPort_6_6;
  assign bankToPort_6_6 = T2506;
  assign T2506 = T2510 ? readValueBankFifo : T2507;
  assign T2507 = T2508 ? readValueBankFifo : 32'h0;
  assign T2508 = T430 & T2509;
  assign T2509 = T1651[3'h6:3'h6];
  assign T2510 = T433 & T2509;
  assign T2511 = T2518 | T2512;
  assign T2512 = bankToPort_5_6;
  assign bankToPort_5_6 = T2513;
  assign T2513 = T2517 ? readValueBankFifo : T2514;
  assign T2514 = T2515 ? readValueBankFifo : 32'h0;
  assign T2515 = T425 & T2516;
  assign T2516 = T1660[3'h6:3'h6];
  assign T2517 = T428 & T2516;
  assign T2518 = T2525 | T2519;
  assign T2519 = bankToPort_4_6;
  assign bankToPort_4_6 = T2520;
  assign T2520 = T2524 ? readValueBankFifo : T2521;
  assign T2521 = T2522 ? readValueBankFifo : 32'h0;
  assign T2522 = T420 & T2523;
  assign T2523 = T1669[3'h6:3'h6];
  assign T2524 = T423 & T2523;
  assign T2525 = T2532 | T2526;
  assign T2526 = bankToPort_3_6;
  assign bankToPort_3_6 = T2527;
  assign T2527 = T2531 ? readValueBankFifo : T2528;
  assign T2528 = T2529 ? readValueBankFifo : 32'h0;
  assign T2529 = T415 & T2530;
  assign T2530 = T1678[3'h6:3'h6];
  assign T2531 = T418 & T2530;
  assign T2532 = T2539 | T2533;
  assign T2533 = bankToPort_2_6;
  assign bankToPort_2_6 = T2534;
  assign T2534 = T2538 ? readValueBankFifo : T2535;
  assign T2535 = T2536 ? readValueBankFifo : 32'h0;
  assign T2536 = T410 & T2537;
  assign T2537 = T1687[3'h6:3'h6];
  assign T2538 = T413 & T2537;
  assign T2539 = T2546 | T2540;
  assign T2540 = bankToPort_1_6;
  assign bankToPort_1_6 = T2541;
  assign T2541 = T2545 ? readValueBankFifo : T2542;
  assign T2542 = T2543 ? readValueBankFifo : 32'h0;
  assign T2543 = T405 & T2544;
  assign T2544 = T1696[3'h6:3'h6];
  assign T2545 = T408 & T2544;
  assign T2546 = 32'h1 | T2547;
  assign T2547 = bankToPort_0_6;
  assign bankToPort_0_6 = T2548;
  assign T2548 = T2552 ? readValueBankFifo : T2549;
  assign T2549 = T2550 ? readValueBankFifo : 32'h0;
  assign T2550 = T402 & T2551;
  assign T2551 = T1705[3'h6:3'h6];
  assign T2552 = T500 & T2551;
  assign T2553 = T781 ^ 1'h1;
  assign T2554 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2555 = T2556 ? 1'h1 : 1'h0;
  assign T2556 = T725 & fifo_25_io_enqRdy;
  assign T2557 = seqLevelDoneReg2 ? fifo_5_io_enqRdy : 1'h0;
  assign T2558 = T2556 ? T2559 : T2559;
  assign T2559 = T2560;
  assign T2560 = T2618 ? 32'h0 : T2561;
  assign T2561 = T725 ? T2562 : 32'h0;
  assign T2562 = T2569 | T2563;
  assign T2563 = bankToPort_7_5;
  assign bankToPort_7_5 = T2564;
  assign T2564 = T2568 ? readValueBankFifo : T2565;
  assign T2565 = T2566 ? readValueBankFifo : 32'h0;
  assign T2566 = T269 & T2567;
  assign T2567 = T1627[3'h5:3'h5];
  assign T2568 = T436 & T2567;
  assign T2569 = T2576 | T2570;
  assign T2570 = bankToPort_6_5;
  assign bankToPort_6_5 = T2571;
  assign T2571 = T2575 ? readValueBankFifo : T2572;
  assign T2572 = T2573 ? readValueBankFifo : 32'h0;
  assign T2573 = T430 & T2574;
  assign T2574 = T1651[3'h5:3'h5];
  assign T2575 = T433 & T2574;
  assign T2576 = T2583 | T2577;
  assign T2577 = bankToPort_5_5;
  assign bankToPort_5_5 = T2578;
  assign T2578 = T2582 ? readValueBankFifo : T2579;
  assign T2579 = T2580 ? readValueBankFifo : 32'h0;
  assign T2580 = T425 & T2581;
  assign T2581 = T1660[3'h5:3'h5];
  assign T2582 = T428 & T2581;
  assign T2583 = T2590 | T2584;
  assign T2584 = bankToPort_4_5;
  assign bankToPort_4_5 = T2585;
  assign T2585 = T2589 ? readValueBankFifo : T2586;
  assign T2586 = T2587 ? readValueBankFifo : 32'h0;
  assign T2587 = T420 & T2588;
  assign T2588 = T1669[3'h5:3'h5];
  assign T2589 = T423 & T2588;
  assign T2590 = T2597 | T2591;
  assign T2591 = bankToPort_3_5;
  assign bankToPort_3_5 = T2592;
  assign T2592 = T2596 ? readValueBankFifo : T2593;
  assign T2593 = T2594 ? readValueBankFifo : 32'h0;
  assign T2594 = T415 & T2595;
  assign T2595 = T1678[3'h5:3'h5];
  assign T2596 = T418 & T2595;
  assign T2597 = T2604 | T2598;
  assign T2598 = bankToPort_2_5;
  assign bankToPort_2_5 = T2599;
  assign T2599 = T2603 ? readValueBankFifo : T2600;
  assign T2600 = T2601 ? readValueBankFifo : 32'h0;
  assign T2601 = T410 & T2602;
  assign T2602 = T1687[3'h5:3'h5];
  assign T2603 = T413 & T2602;
  assign T2604 = T2611 | T2605;
  assign T2605 = bankToPort_1_5;
  assign bankToPort_1_5 = T2606;
  assign T2606 = T2610 ? readValueBankFifo : T2607;
  assign T2607 = T2608 ? readValueBankFifo : 32'h0;
  assign T2608 = T405 & T2609;
  assign T2609 = T1696[3'h5:3'h5];
  assign T2610 = T408 & T2609;
  assign T2611 = 32'h1 | T2612;
  assign T2612 = bankToPort_0_5;
  assign bankToPort_0_5 = T2613;
  assign T2613 = T2617 ? readValueBankFifo : T2614;
  assign T2614 = T2615 ? readValueBankFifo : 32'h0;
  assign T2615 = T402 & T2616;
  assign T2616 = T1705[3'h5:3'h5];
  assign T2617 = T500 & T2616;
  assign T2618 = T725 ^ 1'h1;
  assign T2619 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2620 = T2621 ? 1'h1 : 1'h0;
  assign T2621 = T669 & fifo_24_io_enqRdy;
  assign T2622 = seqLevelDoneReg2 ? fifo_4_io_enqRdy : 1'h0;
  assign T2623 = T2621 ? T2624 : T2624;
  assign T2624 = T2625;
  assign T2625 = T2683 ? 32'h0 : T2626;
  assign T2626 = T669 ? T2627 : 32'h0;
  assign T2627 = T2634 | T2628;
  assign T2628 = bankToPort_7_4;
  assign bankToPort_7_4 = T2629;
  assign T2629 = T2633 ? readValueBankFifo : T2630;
  assign T2630 = T2631 ? readValueBankFifo : 32'h0;
  assign T2631 = T269 & T2632;
  assign T2632 = T1627[3'h4:3'h4];
  assign T2633 = T436 & T2632;
  assign T2634 = T2641 | T2635;
  assign T2635 = bankToPort_6_4;
  assign bankToPort_6_4 = T2636;
  assign T2636 = T2640 ? readValueBankFifo : T2637;
  assign T2637 = T2638 ? readValueBankFifo : 32'h0;
  assign T2638 = T430 & T2639;
  assign T2639 = T1651[3'h4:3'h4];
  assign T2640 = T433 & T2639;
  assign T2641 = T2648 | T2642;
  assign T2642 = bankToPort_5_4;
  assign bankToPort_5_4 = T2643;
  assign T2643 = T2647 ? readValueBankFifo : T2644;
  assign T2644 = T2645 ? readValueBankFifo : 32'h0;
  assign T2645 = T425 & T2646;
  assign T2646 = T1660[3'h4:3'h4];
  assign T2647 = T428 & T2646;
  assign T2648 = T2655 | T2649;
  assign T2649 = bankToPort_4_4;
  assign bankToPort_4_4 = T2650;
  assign T2650 = T2654 ? readValueBankFifo : T2651;
  assign T2651 = T2652 ? readValueBankFifo : 32'h0;
  assign T2652 = T420 & T2653;
  assign T2653 = T1669[3'h4:3'h4];
  assign T2654 = T423 & T2653;
  assign T2655 = T2662 | T2656;
  assign T2656 = bankToPort_3_4;
  assign bankToPort_3_4 = T2657;
  assign T2657 = T2661 ? readValueBankFifo : T2658;
  assign T2658 = T2659 ? readValueBankFifo : 32'h0;
  assign T2659 = T415 & T2660;
  assign T2660 = T1678[3'h4:3'h4];
  assign T2661 = T418 & T2660;
  assign T2662 = T2669 | T2663;
  assign T2663 = bankToPort_2_4;
  assign bankToPort_2_4 = T2664;
  assign T2664 = T2668 ? readValueBankFifo : T2665;
  assign T2665 = T2666 ? readValueBankFifo : 32'h0;
  assign T2666 = T410 & T2667;
  assign T2667 = T1687[3'h4:3'h4];
  assign T2668 = T413 & T2667;
  assign T2669 = T2676 | T2670;
  assign T2670 = bankToPort_1_4;
  assign bankToPort_1_4 = T2671;
  assign T2671 = T2675 ? readValueBankFifo : T2672;
  assign T2672 = T2673 ? readValueBankFifo : 32'h0;
  assign T2673 = T405 & T2674;
  assign T2674 = T1696[3'h4:3'h4];
  assign T2675 = T408 & T2674;
  assign T2676 = 32'h1 | T2677;
  assign T2677 = bankToPort_0_4;
  assign bankToPort_0_4 = T2678;
  assign T2678 = T2682 ? readValueBankFifo : T2679;
  assign T2679 = T2680 ? readValueBankFifo : 32'h0;
  assign T2680 = T402 & T2681;
  assign T2681 = T1705[3'h4:3'h4];
  assign T2682 = T500 & T2681;
  assign T2683 = T669 ^ 1'h1;
  assign T2684 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2685 = T2686 ? 1'h1 : 1'h0;
  assign T2686 = T613 & fifo_23_io_enqRdy;
  assign T2687 = seqLevelDoneReg2 ? fifo_3_io_enqRdy : 1'h0;
  assign T2688 = T2686 ? T2689 : T2689;
  assign T2689 = T2690;
  assign T2690 = T2748 ? 32'h0 : T2691;
  assign T2691 = T613 ? T2692 : 32'h0;
  assign T2692 = T2699 | T2693;
  assign T2693 = bankToPort_7_3;
  assign bankToPort_7_3 = T2694;
  assign T2694 = T2698 ? readValueBankFifo : T2695;
  assign T2695 = T2696 ? readValueBankFifo : 32'h0;
  assign T2696 = T269 & T2697;
  assign T2697 = T1627[2'h3:2'h3];
  assign T2698 = T436 & T2697;
  assign T2699 = T2706 | T2700;
  assign T2700 = bankToPort_6_3;
  assign bankToPort_6_3 = T2701;
  assign T2701 = T2705 ? readValueBankFifo : T2702;
  assign T2702 = T2703 ? readValueBankFifo : 32'h0;
  assign T2703 = T430 & T2704;
  assign T2704 = T1651[2'h3:2'h3];
  assign T2705 = T433 & T2704;
  assign T2706 = T2713 | T2707;
  assign T2707 = bankToPort_5_3;
  assign bankToPort_5_3 = T2708;
  assign T2708 = T2712 ? readValueBankFifo : T2709;
  assign T2709 = T2710 ? readValueBankFifo : 32'h0;
  assign T2710 = T425 & T2711;
  assign T2711 = T1660[2'h3:2'h3];
  assign T2712 = T428 & T2711;
  assign T2713 = T2720 | T2714;
  assign T2714 = bankToPort_4_3;
  assign bankToPort_4_3 = T2715;
  assign T2715 = T2719 ? readValueBankFifo : T2716;
  assign T2716 = T2717 ? readValueBankFifo : 32'h0;
  assign T2717 = T420 & T2718;
  assign T2718 = T1669[2'h3:2'h3];
  assign T2719 = T423 & T2718;
  assign T2720 = T2727 | T2721;
  assign T2721 = bankToPort_3_3;
  assign bankToPort_3_3 = T2722;
  assign T2722 = T2726 ? readValueBankFifo : T2723;
  assign T2723 = T2724 ? readValueBankFifo : 32'h0;
  assign T2724 = T415 & T2725;
  assign T2725 = T1678[2'h3:2'h3];
  assign T2726 = T418 & T2725;
  assign T2727 = T2734 | T2728;
  assign T2728 = bankToPort_2_3;
  assign bankToPort_2_3 = T2729;
  assign T2729 = T2733 ? readValueBankFifo : T2730;
  assign T2730 = T2731 ? readValueBankFifo : 32'h0;
  assign T2731 = T410 & T2732;
  assign T2732 = T1687[2'h3:2'h3];
  assign T2733 = T413 & T2732;
  assign T2734 = T2741 | T2735;
  assign T2735 = bankToPort_1_3;
  assign bankToPort_1_3 = T2736;
  assign T2736 = T2740 ? readValueBankFifo : T2737;
  assign T2737 = T2738 ? readValueBankFifo : 32'h0;
  assign T2738 = T405 & T2739;
  assign T2739 = T1696[2'h3:2'h3];
  assign T2740 = T408 & T2739;
  assign T2741 = 32'h1 | T2742;
  assign T2742 = bankToPort_0_3;
  assign bankToPort_0_3 = T2743;
  assign T2743 = T2747 ? readValueBankFifo : T2744;
  assign T2744 = T2745 ? readValueBankFifo : 32'h0;
  assign T2745 = T402 & T2746;
  assign T2746 = T1705[2'h3:2'h3];
  assign T2747 = T500 & T2746;
  assign T2748 = T613 ^ 1'h1;
  assign T2749 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2750 = T2751 ? 1'h1 : 1'h0;
  assign T2751 = T557 & fifo_22_io_enqRdy;
  assign T2752 = seqLevelDoneReg2 ? fifo_2_io_enqRdy : 1'h0;
  assign T2753 = T2751 ? T2754 : T2754;
  assign T2754 = T2755;
  assign T2755 = T2813 ? 32'h0 : T2756;
  assign T2756 = T557 ? T2757 : 32'h0;
  assign T2757 = T2764 | T2758;
  assign T2758 = bankToPort_7_2;
  assign bankToPort_7_2 = T2759;
  assign T2759 = T2763 ? readValueBankFifo : T2760;
  assign T2760 = T2761 ? readValueBankFifo : 32'h0;
  assign T2761 = T269 & T2762;
  assign T2762 = T1627[2'h2:2'h2];
  assign T2763 = T436 & T2762;
  assign T2764 = T2771 | T2765;
  assign T2765 = bankToPort_6_2;
  assign bankToPort_6_2 = T2766;
  assign T2766 = T2770 ? readValueBankFifo : T2767;
  assign T2767 = T2768 ? readValueBankFifo : 32'h0;
  assign T2768 = T430 & T2769;
  assign T2769 = T1651[2'h2:2'h2];
  assign T2770 = T433 & T2769;
  assign T2771 = T2778 | T2772;
  assign T2772 = bankToPort_5_2;
  assign bankToPort_5_2 = T2773;
  assign T2773 = T2777 ? readValueBankFifo : T2774;
  assign T2774 = T2775 ? readValueBankFifo : 32'h0;
  assign T2775 = T425 & T2776;
  assign T2776 = T1660[2'h2:2'h2];
  assign T2777 = T428 & T2776;
  assign T2778 = T2785 | T2779;
  assign T2779 = bankToPort_4_2;
  assign bankToPort_4_2 = T2780;
  assign T2780 = T2784 ? readValueBankFifo : T2781;
  assign T2781 = T2782 ? readValueBankFifo : 32'h0;
  assign T2782 = T420 & T2783;
  assign T2783 = T1669[2'h2:2'h2];
  assign T2784 = T423 & T2783;
  assign T2785 = T2792 | T2786;
  assign T2786 = bankToPort_3_2;
  assign bankToPort_3_2 = T2787;
  assign T2787 = T2791 ? readValueBankFifo : T2788;
  assign T2788 = T2789 ? readValueBankFifo : 32'h0;
  assign T2789 = T415 & T2790;
  assign T2790 = T1678[2'h2:2'h2];
  assign T2791 = T418 & T2790;
  assign T2792 = T2799 | T2793;
  assign T2793 = bankToPort_2_2;
  assign bankToPort_2_2 = T2794;
  assign T2794 = T2798 ? readValueBankFifo : T2795;
  assign T2795 = T2796 ? readValueBankFifo : 32'h0;
  assign T2796 = T410 & T2797;
  assign T2797 = T1687[2'h2:2'h2];
  assign T2798 = T413 & T2797;
  assign T2799 = T2806 | T2800;
  assign T2800 = bankToPort_1_2;
  assign bankToPort_1_2 = T2801;
  assign T2801 = T2805 ? readValueBankFifo : T2802;
  assign T2802 = T2803 ? readValueBankFifo : 32'h0;
  assign T2803 = T405 & T2804;
  assign T2804 = T1696[2'h2:2'h2];
  assign T2805 = T408 & T2804;
  assign T2806 = 32'h1 | T2807;
  assign T2807 = bankToPort_0_2;
  assign bankToPort_0_2 = T2808;
  assign T2808 = T2812 ? readValueBankFifo : T2809;
  assign T2809 = T2810 ? readValueBankFifo : 32'h0;
  assign T2810 = T402 & T2811;
  assign T2811 = T1705[2'h2:2'h2];
  assign T2812 = T500 & T2811;
  assign T2813 = T557 ^ 1'h1;
  assign T2814 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2815 = T2816 ? 1'h1 : 1'h0;
  assign T2816 = T501 & fifo_21_io_enqRdy;
  assign T2817 = seqLevelDoneReg2 ? fifo_1_io_enqRdy : 1'h0;
  assign T2818 = T2816 ? T2819 : T2819;
  assign T2819 = T2820;
  assign T2820 = T2878 ? 32'h0 : T2821;
  assign T2821 = T501 ? T2822 : 32'h0;
  assign T2822 = T2829 | T2823;
  assign T2823 = bankToPort_7_1;
  assign bankToPort_7_1 = T2824;
  assign T2824 = T2828 ? readValueBankFifo : T2825;
  assign T2825 = T2826 ? readValueBankFifo : 32'h0;
  assign T2826 = T269 & T2827;
  assign T2827 = T1627[1'h1:1'h1];
  assign T2828 = T436 & T2827;
  assign T2829 = T2836 | T2830;
  assign T2830 = bankToPort_6_1;
  assign bankToPort_6_1 = T2831;
  assign T2831 = T2835 ? readValueBankFifo : T2832;
  assign T2832 = T2833 ? readValueBankFifo : 32'h0;
  assign T2833 = T430 & T2834;
  assign T2834 = T1651[1'h1:1'h1];
  assign T2835 = T433 & T2834;
  assign T2836 = T2843 | T2837;
  assign T2837 = bankToPort_5_1;
  assign bankToPort_5_1 = T2838;
  assign T2838 = T2842 ? readValueBankFifo : T2839;
  assign T2839 = T2840 ? readValueBankFifo : 32'h0;
  assign T2840 = T425 & T2841;
  assign T2841 = T1660[1'h1:1'h1];
  assign T2842 = T428 & T2841;
  assign T2843 = T2850 | T2844;
  assign T2844 = bankToPort_4_1;
  assign bankToPort_4_1 = T2845;
  assign T2845 = T2849 ? readValueBankFifo : T2846;
  assign T2846 = T2847 ? readValueBankFifo : 32'h0;
  assign T2847 = T420 & T2848;
  assign T2848 = T1669[1'h1:1'h1];
  assign T2849 = T423 & T2848;
  assign T2850 = T2857 | T2851;
  assign T2851 = bankToPort_3_1;
  assign bankToPort_3_1 = T2852;
  assign T2852 = T2856 ? readValueBankFifo : T2853;
  assign T2853 = T2854 ? readValueBankFifo : 32'h0;
  assign T2854 = T415 & T2855;
  assign T2855 = T1678[1'h1:1'h1];
  assign T2856 = T418 & T2855;
  assign T2857 = T2864 | T2858;
  assign T2858 = bankToPort_2_1;
  assign bankToPort_2_1 = T2859;
  assign T2859 = T2863 ? readValueBankFifo : T2860;
  assign T2860 = T2861 ? readValueBankFifo : 32'h0;
  assign T2861 = T410 & T2862;
  assign T2862 = T1687[1'h1:1'h1];
  assign T2863 = T413 & T2862;
  assign T2864 = T2871 | T2865;
  assign T2865 = bankToPort_1_1;
  assign bankToPort_1_1 = T2866;
  assign T2866 = T2870 ? readValueBankFifo : T2867;
  assign T2867 = T2868 ? readValueBankFifo : 32'h0;
  assign T2868 = T405 & T2869;
  assign T2869 = T1696[1'h1:1'h1];
  assign T2870 = T408 & T2869;
  assign T2871 = 32'h1 | T2872;
  assign T2872 = bankToPort_0_1;
  assign bankToPort_0_1 = T2873;
  assign T2873 = T2877 ? readValueBankFifo : T2874;
  assign T2874 = T2875 ? readValueBankFifo : 32'h0;
  assign T2875 = T402 & T2876;
  assign T2876 = T1705[1'h1:1'h1];
  assign T2877 = T500 & T2876;
  assign T2878 = T501 ^ 1'h1;
  assign T2879 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2880 = T2881 ? 1'h1 : 1'h0;
  assign T2881 = T361 & fifo_20_io_enqRdy;
  assign T2882 = seqLevelDoneReg2 ? fifo_io_enqRdy : 1'h0;
  assign T2883 = T2881 ? T2884 : T2884;
  assign T2884 = T2885;
  assign T2885 = T2943 ? 32'h0 : T2886;
  assign T2886 = T361 ? T2887 : 32'h0;
  assign T2887 = T2894 | T2888;
  assign T2888 = bankToPort_7_0;
  assign bankToPort_7_0 = T2889;
  assign T2889 = T2893 ? readValueBankFifo : T2890;
  assign T2890 = T2891 ? readValueBankFifo : 32'h0;
  assign T2891 = T269 & T2892;
  assign T2892 = T1627[1'h0:1'h0];
  assign T2893 = T436 & T2892;
  assign T2894 = T2901 | T2895;
  assign T2895 = bankToPort_6_0;
  assign bankToPort_6_0 = T2896;
  assign T2896 = T2900 ? readValueBankFifo : T2897;
  assign T2897 = T2898 ? readValueBankFifo : 32'h0;
  assign T2898 = T430 & T2899;
  assign T2899 = T1651[1'h0:1'h0];
  assign T2900 = T433 & T2899;
  assign T2901 = T2908 | T2902;
  assign T2902 = bankToPort_5_0;
  assign bankToPort_5_0 = T2903;
  assign T2903 = T2907 ? readValueBankFifo : T2904;
  assign T2904 = T2905 ? readValueBankFifo : 32'h0;
  assign T2905 = T425 & T2906;
  assign T2906 = T1660[1'h0:1'h0];
  assign T2907 = T428 & T2906;
  assign T2908 = T2915 | T2909;
  assign T2909 = bankToPort_4_0;
  assign bankToPort_4_0 = T2910;
  assign T2910 = T2914 ? readValueBankFifo : T2911;
  assign T2911 = T2912 ? readValueBankFifo : 32'h0;
  assign T2912 = T420 & T2913;
  assign T2913 = T1669[1'h0:1'h0];
  assign T2914 = T423 & T2913;
  assign T2915 = T2922 | T2916;
  assign T2916 = bankToPort_3_0;
  assign bankToPort_3_0 = T2917;
  assign T2917 = T2921 ? readValueBankFifo : T2918;
  assign T2918 = T2919 ? readValueBankFifo : 32'h0;
  assign T2919 = T415 & T2920;
  assign T2920 = T1678[1'h0:1'h0];
  assign T2921 = T418 & T2920;
  assign T2922 = T2929 | T2923;
  assign T2923 = bankToPort_2_0;
  assign bankToPort_2_0 = T2924;
  assign T2924 = T2928 ? readValueBankFifo : T2925;
  assign T2925 = T2926 ? readValueBankFifo : 32'h0;
  assign T2926 = T410 & T2927;
  assign T2927 = T1687[1'h0:1'h0];
  assign T2928 = T413 & T2927;
  assign T2929 = T2936 | T2930;
  assign T2930 = bankToPort_1_0;
  assign bankToPort_1_0 = T2931;
  assign T2931 = T2935 ? readValueBankFifo : T2932;
  assign T2932 = T2933 ? readValueBankFifo : 32'h0;
  assign T2933 = T405 & T2934;
  assign T2934 = T1696[1'h0:1'h0];
  assign T2935 = T408 & T2934;
  assign T2936 = 32'h1 | T2937;
  assign T2937 = bankToPort_0_0;
  assign bankToPort_0_0 = T2938;
  assign T2938 = T2942 ? readValueBankFifo : T2939;
  assign T2939 = T2940 ? readValueBankFifo : 32'h0;
  assign T2940 = T402 & T2941;
  assign T2941 = T1705[1'h0:1'h0];
  assign T2942 = T500 & T2941;
  assign T2943 = T361 ^ 1'h1;
  assign T2944 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2945 = seqLevelDoneReg2 ? fifo_39_io_deqValid : 1'h0;
  assign T2946 = seqLevelDoneReg2 ? fifo_39_io_deqData : fifo_39_io_deqData;
  assign T2947 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2948 = seqLevelDoneReg2 ? fifo_38_io_deqValid : 1'h0;
  assign T2949 = seqLevelDoneReg2 ? fifo_38_io_deqData : fifo_38_io_deqData;
  assign T2950 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2951 = seqLevelDoneReg2 ? fifo_37_io_deqValid : 1'h0;
  assign T2952 = seqLevelDoneReg2 ? fifo_37_io_deqData : fifo_37_io_deqData;
  assign T2953 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2954 = seqLevelDoneReg2 ? fifo_36_io_deqValid : 1'h0;
  assign T2955 = seqLevelDoneReg2 ? fifo_36_io_deqData : fifo_36_io_deqData;
  assign T2956 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2957 = seqLevelDoneReg2 ? fifo_35_io_deqValid : 1'h0;
  assign T2958 = seqLevelDoneReg2 ? fifo_35_io_deqData : fifo_35_io_deqData;
  assign T2959 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2960 = seqLevelDoneReg2 ? fifo_34_io_deqValid : 1'h0;
  assign T2961 = seqLevelDoneReg2 ? fifo_34_io_deqData : fifo_34_io_deqData;
  assign T2962 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2963 = seqLevelDoneReg2 ? fifo_33_io_deqValid : 1'h0;
  assign T2964 = seqLevelDoneReg2 ? fifo_33_io_deqData : fifo_33_io_deqData;
  assign T2965 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2966 = seqLevelDoneReg2 ? fifo_32_io_deqValid : 1'h0;
  assign T2967 = seqLevelDoneReg2 ? fifo_32_io_deqData : fifo_32_io_deqData;
  assign T2968 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2969 = seqLevelDoneReg2 ? fifo_31_io_deqValid : 1'h0;
  assign T2970 = seqLevelDoneReg2 ? fifo_31_io_deqData : fifo_31_io_deqData;
  assign T2971 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2972 = seqLevelDoneReg2 ? fifo_30_io_deqValid : 1'h0;
  assign T2973 = seqLevelDoneReg2 ? fifo_30_io_deqData : fifo_30_io_deqData;
  assign T2974 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2975 = seqLevelDoneReg2 ? fifo_29_io_deqValid : 1'h0;
  assign T2976 = seqLevelDoneReg2 ? fifo_29_io_deqData : fifo_29_io_deqData;
  assign T2977 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2978 = seqLevelDoneReg2 ? fifo_28_io_deqValid : 1'h0;
  assign T2979 = seqLevelDoneReg2 ? fifo_28_io_deqData : fifo_28_io_deqData;
  assign T2980 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2981 = seqLevelDoneReg2 ? fifo_27_io_deqValid : 1'h0;
  assign T2982 = seqLevelDoneReg2 ? fifo_27_io_deqData : fifo_27_io_deqData;
  assign T2983 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2984 = seqLevelDoneReg2 ? fifo_26_io_deqValid : 1'h0;
  assign T2985 = seqLevelDoneReg2 ? fifo_26_io_deqData : fifo_26_io_deqData;
  assign T2986 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2987 = seqLevelDoneReg2 ? fifo_25_io_deqValid : 1'h0;
  assign T2988 = seqLevelDoneReg2 ? fifo_25_io_deqData : fifo_25_io_deqData;
  assign T2989 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2990 = seqLevelDoneReg2 ? fifo_24_io_deqValid : 1'h0;
  assign T2991 = seqLevelDoneReg2 ? fifo_24_io_deqData : fifo_24_io_deqData;
  assign T2992 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2993 = seqLevelDoneReg2 ? fifo_23_io_deqValid : 1'h0;
  assign T2994 = seqLevelDoneReg2 ? fifo_23_io_deqData : fifo_23_io_deqData;
  assign T2995 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2996 = seqLevelDoneReg2 ? fifo_22_io_deqValid : 1'h0;
  assign T2997 = seqLevelDoneReg2 ? fifo_22_io_deqData : fifo_22_io_deqData;
  assign T2998 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T2999 = seqLevelDoneReg2 ? fifo_21_io_deqValid : 1'h0;
  assign T3000 = seqLevelDoneReg2 ? fifo_21_io_deqData : fifo_21_io_deqData;
  assign T3001 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T3002 = seqLevelDoneReg2 ? fifo_20_io_deqValid : 1'h0;
  assign T3003 = seqLevelDoneReg2 ? fifo_20_io_deqData : fifo_20_io_deqData;
  assign T3004 = fabInSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T3005 = T3009 ? 1'h0 : T3006;
  assign T3006 = T3007 ? 1'h1 : 1'h0;
  assign T3007 = T17 & T3008;
  assign T3008 = bankSeq[7'h56:7'h56];
  assign T3009 = T17 & T3010;
  assign T3010 = T3008 ^ 1'h1;
  assign T3011 = T3015 ? 1'h0 : T3012;
  assign T3012 = T3013 ? 1'h1 : 1'h0;
  assign T3013 = T254 & T3014;
  assign T3014 = bankSeq[7'h56:7'h56];
  assign T3015 = T254 & T3016;
  assign T3016 = T3014 ^ 1'h1;
  assign T3017 = T3021 ? 1'h0 : T3018;
  assign T3018 = T3019 ? 1'h1 : 1'h0;
  assign T3019 = T256 & T3020;
  assign T3020 = bankSeq[7'h56:7'h56];
  assign T3021 = T256 & T3022;
  assign T3022 = T3020 ^ 1'h1;
  assign T3023 = T3027 ? 1'h0 : T3024;
  assign T3024 = T3025 ? 1'h1 : 1'h0;
  assign T3025 = T258 & T3026;
  assign T3026 = bankSeq[7'h56:7'h56];
  assign T3027 = T258 & T3028;
  assign T3028 = T3026 ^ 1'h1;
  assign T3029 = T3033 ? 1'h0 : T3030;
  assign T3030 = T3031 ? 1'h1 : 1'h0;
  assign T3031 = T260 & T3032;
  assign T3032 = bankSeq[7'h56:7'h56];
  assign T3033 = T260 & T3034;
  assign T3034 = T3032 ^ 1'h1;
  assign T3035 = T3039 ? 1'h0 : T3036;
  assign T3036 = T3037 ? 1'h1 : 1'h0;
  assign T3037 = T262 & T3038;
  assign T3038 = bankSeq[7'h56:7'h56];
  assign T3039 = T262 & T3040;
  assign T3040 = T3038 ^ 1'h1;
  assign T3041 = T3045 ? 1'h0 : T3042;
  assign T3042 = T3043 ? 1'h1 : 1'h0;
  assign T3043 = T264 & T3044;
  assign T3044 = bankSeq[7'h56:7'h56];
  assign T3045 = T264 & T3046;
  assign T3046 = T3044 ^ 1'h1;
  assign T3047 = T3051 ? 1'h0 : T3048;
  assign T3048 = T3049 ? 1'h1 : 1'h0;
  assign T3049 = T267 & T3050;
  assign T3050 = bankSeq[7'h56:7'h56];
  assign T3051 = T267 & T3052;
  assign T3052 = T3050 ^ 1'h1;
  assign T3053 = T17 ? 1'h1 : 1'h0;
  assign T3054 = T254 ? 1'h1 : 1'h0;
  assign T3055 = T256 ? 1'h1 : 1'h0;
  assign T3056 = T258 ? 1'h1 : 1'h0;
  assign T3057 = T260 ? 1'h1 : 1'h0;
  assign T3058 = T262 ? 1'h1 : 1'h0;
  assign T3059 = T264 ? 1'h1 : 1'h0;
  assign T3060 = T267 ? 1'h1 : 1'h0;
  assign T3061 = T17 ? readAddr : 6'h0;
  assign readAddr = T3062;
  assign T3062 = T266 ? 6'h0 : T3063;
  assign T3063 = T240 ? T3084 : T3064;
  assign T3064 = T265 ? 6'h0 : T3065;
  assign T3065 = T232 ? T3083 : T3066;
  assign T3066 = T263 ? 6'h0 : T3067;
  assign T3067 = T224 ? T3082 : T3068;
  assign T3068 = T261 ? 6'h0 : T3069;
  assign T3069 = T216 ? T3081 : T3070;
  assign T3070 = T259 ? 6'h0 : T3071;
  assign T3071 = T208 ? T3080 : T3072;
  assign T3072 = T257 ? 6'h0 : T3073;
  assign T3073 = T200 ? T3079 : T3074;
  assign T3074 = T255 ? 6'h0 : T3075;
  assign T3075 = T183 ? T3078 : T3076;
  assign T3076 = T247 ? T3077 : 6'h0;
  assign T3077 = bankSeq[4'h8:2'h3];
  assign T3078 = bankSeq[4'h8:2'h3];
  assign T3079 = bankSeq[4'h8:2'h3];
  assign T3080 = bankSeq[4'h8:2'h3];
  assign T3081 = bankSeq[4'h8:2'h3];
  assign T3082 = bankSeq[4'h8:2'h3];
  assign T3083 = bankSeq[4'h8:2'h3];
  assign T3084 = bankSeq[4'h8:2'h3];
  assign T3085 = T254 ? readAddr : 6'h0;
  assign T3086 = T256 ? readAddr : 6'h0;
  assign T3087 = T258 ? readAddr : 6'h0;
  assign T3088 = T260 ? readAddr : 6'h0;
  assign T3089 = T262 ? readAddr : 6'h0;
  assign T3090 = T264 ? readAddr : 6'h0;
  assign T3091 = T267 ? readAddr : 6'h0;
  assign T3092 = io_seqMemAddrValid ? io_seqMemAddr : io_seqMemAddr;
  assign T3093 = io_seqMemAddrValid ? io_seqMemAddrValid : io_seqMemAddrValid;
  assign io_seqProceed = T3094;
  assign T3094 = T3095 ? 1'h1 : 1'h0;
  assign T3095 = T3097 | T3096;
  assign T3096 = ~ nextSeqRegValid2;
  assign T3097 = ~ nextSeqRegValid1;
  assign io_fabStoreRdy_0 = localStorage_io_enqRdyFabric_0;
  assign io_fabStoreRdy_1 = localStorage_io_enqRdyFabric_1;
  assign io_fabStoreRdy_2 = localStorage_io_enqRdyFabric_2;
  assign io_fabStoreRdy_3 = localStorage_io_enqRdyFabric_3;
  assign io_fabStoreRdy_4 = localStorage_io_enqRdyFabric_4;
  assign io_fabStoreRdy_5 = localStorage_io_enqRdyFabric_5;
  assign io_fabStoreRdy_6 = localStorage_io_enqRdyFabric_6;
  assign io_fabStoreRdy_7 = localStorage_io_enqRdyFabric_7;
  assign io_loadStoreRdy_0 = localStorage_io_enqRdyLoad_0;
  assign io_loadStoreRdy_1 = localStorage_io_enqRdyLoad_1;
  assign io_loadStoreRdy_2 = localStorage_io_enqRdyLoad_2;
  assign io_loadStoreRdy_3 = localStorage_io_enqRdyLoad_3;
  assign io_loadStoreRdy_4 = localStorage_io_enqRdyLoad_4;
  assign io_loadStoreRdy_5 = localStorage_io_enqRdyLoad_5;
  assign io_loadStoreRdy_6 = localStorage_io_enqRdyLoad_6;
  assign io_loadStoreRdy_7 = localStorage_io_enqRdyLoad_7;
  assign io_fabInValid_0 = fifo_io_deqValid;
  assign io_fabInValid_1 = fifo_1_io_deqValid;
  assign io_fabInValid_2 = fifo_2_io_deqValid;
  assign io_fabInValid_3 = fifo_3_io_deqValid;
  assign io_fabInValid_4 = fifo_4_io_deqValid;
  assign io_fabInValid_5 = fifo_5_io_deqValid;
  assign io_fabInValid_6 = fifo_6_io_deqValid;
  assign io_fabInValid_7 = fifo_7_io_deqValid;
  assign io_fabInValid_8 = fifo_8_io_deqValid;
  assign io_fabInValid_9 = fifo_9_io_deqValid;
  assign io_fabInValid_10 = fifo_10_io_deqValid;
  assign io_fabInValid_11 = fifo_11_io_deqValid;
  assign io_fabInValid_12 = fifo_12_io_deqValid;
  assign io_fabInValid_13 = fifo_13_io_deqValid;
  assign io_fabInValid_14 = fifo_14_io_deqValid;
  assign io_fabInValid_15 = fifo_15_io_deqValid;
  assign io_fabInValid_16 = fifo_16_io_deqValid;
  assign io_fabInValid_17 = fifo_17_io_deqValid;
  assign io_fabInValid_18 = fifo_18_io_deqValid;
  assign io_fabInValid_19 = fifo_19_io_deqValid;
  assign io_fabInData_0 = fifo_io_deqData;
  assign io_fabInData_1 = fifo_1_io_deqData;
  assign io_fabInData_2 = fifo_2_io_deqData;
  assign io_fabInData_3 = fifo_3_io_deqData;
  assign io_fabInData_4 = fifo_4_io_deqData;
  assign io_fabInData_5 = fifo_5_io_deqData;
  assign io_fabInData_6 = fifo_6_io_deqData;
  assign io_fabInData_7 = fifo_7_io_deqData;
  assign io_fabInData_8 = fifo_8_io_deqData;
  assign io_fabInData_9 = fifo_9_io_deqData;
  assign io_fabInData_10 = fifo_10_io_deqData;
  assign io_fabInData_11 = fifo_11_io_deqData;
  assign io_fabInData_12 = fifo_12_io_deqData;
  assign io_fabInData_13 = fifo_13_io_deqData;
  assign io_fabInData_14 = fifo_14_io_deqData;
  assign io_fabInData_15 = fifo_15_io_deqData;
  assign io_fabInData_16 = fifo_16_io_deqData;
  assign io_fabInData_17 = fifo_17_io_deqData;
  assign io_fabInData_18 = fifo_18_io_deqData;
  assign io_fabInData_19 = fifo_19_io_deqData;
  customReg_0 fabInSeqMem(.clk(clk),
       .io_inData( fabInSeqMemConfig_io_memData ),
       .io_outData( fabInSeqMem_io_outData ),
       .io_readEn( T3093 ),
       .io_writeEn( fabInSeqMemConfig_io_memOutValid ),
       .io_readAddr( T3092 ),
       .io_writeAddr( fabInSeqMemConfig_io_memAddr )
  );
  controllerLocalStorage localStorage(.clk(clk), .reset(reset),
       .io_inDataLoad_7( io_loadStore_7 ),
       .io_inDataLoad_6( io_loadStore_6 ),
       .io_inDataLoad_5( io_loadStore_5 ),
       .io_inDataLoad_4( io_loadStore_4 ),
       .io_inDataLoad_3( io_loadStore_3 ),
       .io_inDataLoad_2( io_loadStore_2 ),
       .io_inDataLoad_1( io_loadStore_1 ),
       .io_inDataLoad_0( io_loadStore_0 ),
       .io_inDataFabric_7( io_fabStore_7 ),
       .io_inDataFabric_6( io_fabStore_6 ),
       .io_inDataFabric_5( io_fabStore_5 ),
       .io_inDataFabric_4( io_fabStore_4 ),
       .io_inDataFabric_3( io_fabStore_3 ),
       .io_inDataFabric_2( io_fabStore_2 ),
       .io_inDataFabric_1( io_fabStore_1 ),
       .io_inDataFabric_0( io_fabStore_0 ),
       .io_outData_7( localStorage_io_outData_7 ),
       .io_outData_6( localStorage_io_outData_6 ),
       .io_outData_5( localStorage_io_outData_5 ),
       .io_outData_4( localStorage_io_outData_4 ),
       .io_outData_3( localStorage_io_outData_3 ),
       .io_outData_2( localStorage_io_outData_2 ),
       .io_outData_1( localStorage_io_outData_1 ),
       .io_outData_0( localStorage_io_outData_0 ),
       .io_isReadValid_7( localStorage_io_isReadValid_7 ),
       .io_isReadValid_6( localStorage_io_isReadValid_6 ),
       .io_isReadValid_5( localStorage_io_isReadValid_5 ),
       .io_isReadValid_4( localStorage_io_isReadValid_4 ),
       .io_isReadValid_3( localStorage_io_isReadValid_3 ),
       .io_isReadValid_2( localStorage_io_isReadValid_2 ),
       .io_isReadValid_1( localStorage_io_isReadValid_1 ),
       .io_isReadValid_0( localStorage_io_isReadValid_0 ),
       .io_readAddr_7( T3091 ),
       .io_readAddr_6( T3090 ),
       .io_readAddr_5( T3089 ),
       .io_readAddr_4( T3088 ),
       .io_readAddr_3( T3087 ),
       .io_readAddr_2( T3086 ),
       .io_readAddr_1( T3085 ),
       .io_readAddr_0( T3061 ),
       .io_readEn_7( T3060 ),
       .io_readEn_6( T3059 ),
       .io_readEn_5( T3058 ),
       .io_readEn_4( T3057 ),
       .io_readEn_3( T3056 ),
       .io_readEn_2( T3055 ),
       .io_readEn_1( T3054 ),
       .io_readEn_0( T3053 ),
       .io_doInvalidate_7( T3047 ),
       .io_doInvalidate_6( T3041 ),
       .io_doInvalidate_5( T3035 ),
       .io_doInvalidate_4( T3029 ),
       .io_doInvalidate_3( T3023 ),
       .io_doInvalidate_2( T3017 ),
       .io_doInvalidate_1( T3011 ),
       .io_doInvalidate_0( T3005 ),
       //.io_readSuccess_7(  )
       //.io_readSuccess_6(  )
       //.io_readSuccess_5(  )
       //.io_readSuccess_4(  )
       //.io_readSuccess_3(  )
       //.io_readSuccess_2(  )
       //.io_readSuccess_1(  )
       //.io_readSuccess_0(  )
       //.io_writeSuccess_7(  )
       //.io_writeSuccess_6(  )
       //.io_writeSuccess_5(  )
       //.io_writeSuccess_4(  )
       //.io_writeSuccess_3(  )
       //.io_writeSuccess_2(  )
       //.io_writeSuccess_1(  )
       //.io_writeSuccess_0(  )
       .io_enqRdyLoad_7( localStorage_io_enqRdyLoad_7 ),
       .io_enqRdyLoad_6( localStorage_io_enqRdyLoad_6 ),
       .io_enqRdyLoad_5( localStorage_io_enqRdyLoad_5 ),
       .io_enqRdyLoad_4( localStorage_io_enqRdyLoad_4 ),
       .io_enqRdyLoad_3( localStorage_io_enqRdyLoad_3 ),
       .io_enqRdyLoad_2( localStorage_io_enqRdyLoad_2 ),
       .io_enqRdyLoad_1( localStorage_io_enqRdyLoad_1 ),
       .io_enqRdyLoad_0( localStorage_io_enqRdyLoad_0 ),
       .io_enqRdyFabric_7( localStorage_io_enqRdyFabric_7 ),
       .io_enqRdyFabric_6( localStorage_io_enqRdyFabric_6 ),
       .io_enqRdyFabric_5( localStorage_io_enqRdyFabric_5 ),
       .io_enqRdyFabric_4( localStorage_io_enqRdyFabric_4 ),
       .io_enqRdyFabric_3( localStorage_io_enqRdyFabric_3 ),
       .io_enqRdyFabric_2( localStorage_io_enqRdyFabric_2 ),
       .io_enqRdyFabric_1( localStorage_io_enqRdyFabric_1 ),
       .io_enqRdyFabric_0( localStorage_io_enqRdyFabric_0 ),
       .io_enqValidLoad_7( io_loadStoreValid_7 ),
       .io_enqValidLoad_6( io_loadStoreValid_6 ),
       .io_enqValidLoad_5( io_loadStoreValid_5 ),
       .io_enqValidLoad_4( io_loadStoreValid_4 ),
       .io_enqValidLoad_3( io_loadStoreValid_3 ),
       .io_enqValidLoad_2( io_loadStoreValid_2 ),
       .io_enqValidLoad_1( io_loadStoreValid_1 ),
       .io_enqValidLoad_0( io_loadStoreValid_0 ),
       .io_enqValidFabric_7( io_fabStoreValid_7 ),
       .io_enqValidFabric_6( io_fabStoreValid_6 ),
       .io_enqValidFabric_5( io_fabStoreValid_5 ),
       .io_enqValidFabric_4( io_fabStoreValid_4 ),
       .io_enqValidFabric_3( io_fabStoreValid_3 ),
       .io_enqValidFabric_2( io_fabStoreValid_2 ),
       .io_enqValidFabric_1( io_fabStoreValid_1 ),
       .io_enqValidFabric_0( io_fabStoreValid_0 ),
       .io_rst( T3004 )
  );
  memConfig_0 fabInSeqMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( fabInSeqMemConfig_io_memAddr ),
       .io_memData( fabInSeqMemConfig_io_memData ),
       .io_memOutValid( fabInSeqMemConfig_io_memOutValid ),
       .io_rst( fabInSeqMemConfig_io_rst )
  );
  fifo_0 fifo(.clk(clk), .reset(reset),
       .io_enqData( T3003 ),
       .io_deqData( fifo_io_deqData ),
       .io_enqRdy( fifo_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_0 ),
       .io_enqValid( T3002 ),
       .io_deqValid( fifo_io_deqValid ),
       .io_rst( T3001 )
  );
  fifo_0 fifo_1(.clk(clk), .reset(reset),
       .io_enqData( T3000 ),
       .io_deqData( fifo_1_io_deqData ),
       .io_enqRdy( fifo_1_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_1 ),
       .io_enqValid( T2999 ),
       .io_deqValid( fifo_1_io_deqValid ),
       .io_rst( T2998 )
  );
  fifo_0 fifo_2(.clk(clk), .reset(reset),
       .io_enqData( T2997 ),
       .io_deqData( fifo_2_io_deqData ),
       .io_enqRdy( fifo_2_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_2 ),
       .io_enqValid( T2996 ),
       .io_deqValid( fifo_2_io_deqValid ),
       .io_rst( T2995 )
  );
  fifo_0 fifo_3(.clk(clk), .reset(reset),
       .io_enqData( T2994 ),
       .io_deqData( fifo_3_io_deqData ),
       .io_enqRdy( fifo_3_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_3 ),
       .io_enqValid( T2993 ),
       .io_deqValid( fifo_3_io_deqValid ),
       .io_rst( T2992 )
  );
  fifo_0 fifo_4(.clk(clk), .reset(reset),
       .io_enqData( T2991 ),
       .io_deqData( fifo_4_io_deqData ),
       .io_enqRdy( fifo_4_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_4 ),
       .io_enqValid( T2990 ),
       .io_deqValid( fifo_4_io_deqValid ),
       .io_rst( T2989 )
  );
  fifo_0 fifo_5(.clk(clk), .reset(reset),
       .io_enqData( T2988 ),
       .io_deqData( fifo_5_io_deqData ),
       .io_enqRdy( fifo_5_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_5 ),
       .io_enqValid( T2987 ),
       .io_deqValid( fifo_5_io_deqValid ),
       .io_rst( T2986 )
  );
  fifo_0 fifo_6(.clk(clk), .reset(reset),
       .io_enqData( T2985 ),
       .io_deqData( fifo_6_io_deqData ),
       .io_enqRdy( fifo_6_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_6 ),
       .io_enqValid( T2984 ),
       .io_deqValid( fifo_6_io_deqValid ),
       .io_rst( T2983 )
  );
  fifo_0 fifo_7(.clk(clk), .reset(reset),
       .io_enqData( T2982 ),
       .io_deqData( fifo_7_io_deqData ),
       .io_enqRdy( fifo_7_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_7 ),
       .io_enqValid( T2981 ),
       .io_deqValid( fifo_7_io_deqValid ),
       .io_rst( T2980 )
  );
  fifo_0 fifo_8(.clk(clk), .reset(reset),
       .io_enqData( T2979 ),
       .io_deqData( fifo_8_io_deqData ),
       .io_enqRdy( fifo_8_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_8 ),
       .io_enqValid( T2978 ),
       .io_deqValid( fifo_8_io_deqValid ),
       .io_rst( T2977 )
  );
  fifo_0 fifo_9(.clk(clk), .reset(reset),
       .io_enqData( T2976 ),
       .io_deqData( fifo_9_io_deqData ),
       .io_enqRdy( fifo_9_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_9 ),
       .io_enqValid( T2975 ),
       .io_deqValid( fifo_9_io_deqValid ),
       .io_rst( T2974 )
  );
  fifo_0 fifo_10(.clk(clk), .reset(reset),
       .io_enqData( T2973 ),
       .io_deqData( fifo_10_io_deqData ),
       .io_enqRdy( fifo_10_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_10 ),
       .io_enqValid( T2972 ),
       .io_deqValid( fifo_10_io_deqValid ),
       .io_rst( T2971 )
  );
  fifo_0 fifo_11(.clk(clk), .reset(reset),
       .io_enqData( T2970 ),
       .io_deqData( fifo_11_io_deqData ),
       .io_enqRdy( fifo_11_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_11 ),
       .io_enqValid( T2969 ),
       .io_deqValid( fifo_11_io_deqValid ),
       .io_rst( T2968 )
  );
  fifo_0 fifo_12(.clk(clk), .reset(reset),
       .io_enqData( T2967 ),
       .io_deqData( fifo_12_io_deqData ),
       .io_enqRdy( fifo_12_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_12 ),
       .io_enqValid( T2966 ),
       .io_deqValid( fifo_12_io_deqValid ),
       .io_rst( T2965 )
  );
  fifo_0 fifo_13(.clk(clk), .reset(reset),
       .io_enqData( T2964 ),
       .io_deqData( fifo_13_io_deqData ),
       .io_enqRdy( fifo_13_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_13 ),
       .io_enqValid( T2963 ),
       .io_deqValid( fifo_13_io_deqValid ),
       .io_rst( T2962 )
  );
  fifo_0 fifo_14(.clk(clk), .reset(reset),
       .io_enqData( T2961 ),
       .io_deqData( fifo_14_io_deqData ),
       .io_enqRdy( fifo_14_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_14 ),
       .io_enqValid( T2960 ),
       .io_deqValid( fifo_14_io_deqValid ),
       .io_rst( T2959 )
  );
  fifo_0 fifo_15(.clk(clk), .reset(reset),
       .io_enqData( T2958 ),
       .io_deqData( fifo_15_io_deqData ),
       .io_enqRdy( fifo_15_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_15 ),
       .io_enqValid( T2957 ),
       .io_deqValid( fifo_15_io_deqValid ),
       .io_rst( T2956 )
  );
  fifo_0 fifo_16(.clk(clk), .reset(reset),
       .io_enqData( T2955 ),
       .io_deqData( fifo_16_io_deqData ),
       .io_enqRdy( fifo_16_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_16 ),
       .io_enqValid( T2954 ),
       .io_deqValid( fifo_16_io_deqValid ),
       .io_rst( T2953 )
  );
  fifo_0 fifo_17(.clk(clk), .reset(reset),
       .io_enqData( T2952 ),
       .io_deqData( fifo_17_io_deqData ),
       .io_enqRdy( fifo_17_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_17 ),
       .io_enqValid( T2951 ),
       .io_deqValid( fifo_17_io_deqValid ),
       .io_rst( T2950 )
  );
  fifo_0 fifo_18(.clk(clk), .reset(reset),
       .io_enqData( T2949 ),
       .io_deqData( fifo_18_io_deqData ),
       .io_enqRdy( fifo_18_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_18 ),
       .io_enqValid( T2948 ),
       .io_deqValid( fifo_18_io_deqValid ),
       .io_rst( T2947 )
  );
  fifo_0 fifo_19(.clk(clk), .reset(reset),
       .io_enqData( T2946 ),
       .io_deqData( fifo_19_io_deqData ),
       .io_enqRdy( fifo_19_io_enqRdy ),
       .io_deqRdy( io_fabInRdy_19 ),
       .io_enqValid( T2945 ),
       .io_deqValid( fifo_19_io_deqValid ),
       .io_rst( T2944 )
  );
  fifo_1 fifo_20(.clk(clk), .reset(reset),
       .io_enqData( T2883 ),
       .io_deqData( fifo_20_io_deqData ),
       .io_enqRdy( fifo_20_io_enqRdy ),
       .io_deqRdy( T2882 ),
       .io_enqValid( T2880 ),
       .io_deqValid( fifo_20_io_deqValid ),
       .io_rst( T2879 )
  );
  fifo_1 fifo_21(.clk(clk), .reset(reset),
       .io_enqData( T2818 ),
       .io_deqData( fifo_21_io_deqData ),
       .io_enqRdy( fifo_21_io_enqRdy ),
       .io_deqRdy( T2817 ),
       .io_enqValid( T2815 ),
       .io_deqValid( fifo_21_io_deqValid ),
       .io_rst( T2814 )
  );
  fifo_1 fifo_22(.clk(clk), .reset(reset),
       .io_enqData( T2753 ),
       .io_deqData( fifo_22_io_deqData ),
       .io_enqRdy( fifo_22_io_enqRdy ),
       .io_deqRdy( T2752 ),
       .io_enqValid( T2750 ),
       .io_deqValid( fifo_22_io_deqValid ),
       .io_rst( T2749 )
  );
  fifo_1 fifo_23(.clk(clk), .reset(reset),
       .io_enqData( T2688 ),
       .io_deqData( fifo_23_io_deqData ),
       .io_enqRdy( fifo_23_io_enqRdy ),
       .io_deqRdy( T2687 ),
       .io_enqValid( T2685 ),
       .io_deqValid( fifo_23_io_deqValid ),
       .io_rst( T2684 )
  );
  fifo_1 fifo_24(.clk(clk), .reset(reset),
       .io_enqData( T2623 ),
       .io_deqData( fifo_24_io_deqData ),
       .io_enqRdy( fifo_24_io_enqRdy ),
       .io_deqRdy( T2622 ),
       .io_enqValid( T2620 ),
       .io_deqValid( fifo_24_io_deqValid ),
       .io_rst( T2619 )
  );
  fifo_1 fifo_25(.clk(clk), .reset(reset),
       .io_enqData( T2558 ),
       .io_deqData( fifo_25_io_deqData ),
       .io_enqRdy( fifo_25_io_enqRdy ),
       .io_deqRdy( T2557 ),
       .io_enqValid( T2555 ),
       .io_deqValid( fifo_25_io_deqValid ),
       .io_rst( T2554 )
  );
  fifo_1 fifo_26(.clk(clk), .reset(reset),
       .io_enqData( T2493 ),
       .io_deqData( fifo_26_io_deqData ),
       .io_enqRdy( fifo_26_io_enqRdy ),
       .io_deqRdy( T2492 ),
       .io_enqValid( T2490 ),
       .io_deqValid( fifo_26_io_deqValid ),
       .io_rst( T2489 )
  );
  fifo_1 fifo_27(.clk(clk), .reset(reset),
       .io_enqData( T2428 ),
       .io_deqData( fifo_27_io_deqData ),
       .io_enqRdy( fifo_27_io_enqRdy ),
       .io_deqRdy( T2427 ),
       .io_enqValid( T2425 ),
       .io_deqValid( fifo_27_io_deqValid ),
       .io_rst( T2424 )
  );
  fifo_1 fifo_28(.clk(clk), .reset(reset),
       .io_enqData( T2363 ),
       .io_deqData( fifo_28_io_deqData ),
       .io_enqRdy( fifo_28_io_enqRdy ),
       .io_deqRdy( T2362 ),
       .io_enqValid( T2360 ),
       .io_deqValid( fifo_28_io_deqValid ),
       .io_rst( T2359 )
  );
  fifo_1 fifo_29(.clk(clk), .reset(reset),
       .io_enqData( T2298 ),
       .io_deqData( fifo_29_io_deqData ),
       .io_enqRdy( fifo_29_io_enqRdy ),
       .io_deqRdy( T2297 ),
       .io_enqValid( T2295 ),
       .io_deqValid( fifo_29_io_deqValid ),
       .io_rst( T2294 )
  );
  fifo_1 fifo_30(.clk(clk), .reset(reset),
       .io_enqData( T2233 ),
       .io_deqData( fifo_30_io_deqData ),
       .io_enqRdy( fifo_30_io_enqRdy ),
       .io_deqRdy( T2232 ),
       .io_enqValid( T2230 ),
       .io_deqValid( fifo_30_io_deqValid ),
       .io_rst( T2229 )
  );
  fifo_1 fifo_31(.clk(clk), .reset(reset),
       .io_enqData( T2168 ),
       .io_deqData( fifo_31_io_deqData ),
       .io_enqRdy( fifo_31_io_enqRdy ),
       .io_deqRdy( T2167 ),
       .io_enqValid( T2165 ),
       .io_deqValid( fifo_31_io_deqValid ),
       .io_rst( T2164 )
  );
  fifo_1 fifo_32(.clk(clk), .reset(reset),
       .io_enqData( T2103 ),
       .io_deqData( fifo_32_io_deqData ),
       .io_enqRdy( fifo_32_io_enqRdy ),
       .io_deqRdy( T2102 ),
       .io_enqValid( T2100 ),
       .io_deqValid( fifo_32_io_deqValid ),
       .io_rst( T2099 )
  );
  fifo_1 fifo_33(.clk(clk), .reset(reset),
       .io_enqData( T2038 ),
       .io_deqData( fifo_33_io_deqData ),
       .io_enqRdy( fifo_33_io_enqRdy ),
       .io_deqRdy( T2037 ),
       .io_enqValid( T2035 ),
       .io_deqValid( fifo_33_io_deqValid ),
       .io_rst( T2034 )
  );
  fifo_1 fifo_34(.clk(clk), .reset(reset),
       .io_enqData( T1973 ),
       .io_deqData( fifo_34_io_deqData ),
       .io_enqRdy( fifo_34_io_enqRdy ),
       .io_deqRdy( T1972 ),
       .io_enqValid( T1970 ),
       .io_deqValid( fifo_34_io_deqValid ),
       .io_rst( T1969 )
  );
  fifo_1 fifo_35(.clk(clk), .reset(reset),
       .io_enqData( T1908 ),
       .io_deqData( fifo_35_io_deqData ),
       .io_enqRdy( fifo_35_io_enqRdy ),
       .io_deqRdy( T1907 ),
       .io_enqValid( T1905 ),
       .io_deqValid( fifo_35_io_deqValid ),
       .io_rst( T1904 )
  );
  fifo_1 fifo_36(.clk(clk), .reset(reset),
       .io_enqData( T1843 ),
       .io_deqData( fifo_36_io_deqData ),
       .io_enqRdy( fifo_36_io_enqRdy ),
       .io_deqRdy( T1842 ),
       .io_enqValid( T1840 ),
       .io_deqValid( fifo_36_io_deqValid ),
       .io_rst( T1839 )
  );
  fifo_1 fifo_37(.clk(clk), .reset(reset),
       .io_enqData( T1778 ),
       .io_deqData( fifo_37_io_deqData ),
       .io_enqRdy( fifo_37_io_enqRdy ),
       .io_deqRdy( T1777 ),
       .io_enqValid( T1775 ),
       .io_deqValid( fifo_37_io_deqValid ),
       .io_rst( T1774 )
  );
  fifo_1 fifo_38(.clk(clk), .reset(reset),
       .io_enqData( T1713 ),
       .io_deqData( fifo_38_io_deqData ),
       .io_enqRdy( fifo_38_io_enqRdy ),
       .io_deqRdy( T1712 ),
       .io_enqValid( T1710 ),
       .io_deqValid( fifo_38_io_deqValid ),
       .io_rst( T1709 )
  );
  fifo_1 fifo_39(.clk(clk), .reset(reset),
       .io_enqData( T1617 ),
       .io_deqData( fifo_39_io_deqData ),
       .io_enqRdy( fifo_39_io_enqRdy ),
       .io_deqRdy( T1616 ),
       .io_enqValid( T1614 ),
       .io_deqValid( fifo_39_io_deqValid ),
       .io_rst( T1613 )
  );
  fifo_0 fifo_40(.clk(clk), .reset(reset),
       .io_enqData( T1612 ),
       .io_deqData( fifo_40_io_deqData ),
       .io_enqRdy( fifo_40_io_enqRdy ),
       .io_deqRdy( T1611 ),
       .io_enqValid( T1610 ),
       .io_deqValid( fifo_40_io_deqValid ),
       .io_rst( T1609 )
  );
  fifo_0 fifo_41(.clk(clk), .reset(reset),
       .io_enqData( T1608 ),
       .io_deqData( fifo_41_io_deqData ),
       .io_enqRdy( fifo_41_io_enqRdy ),
       .io_deqRdy( T1607 ),
       .io_enqValid( T1606 ),
       .io_deqValid( fifo_41_io_deqValid ),
       .io_rst( T1605 )
  );
  fifo_0 fifo_42(.clk(clk), .reset(reset),
       .io_enqData( T1604 ),
       .io_deqData( fifo_42_io_deqData ),
       .io_enqRdy( fifo_42_io_enqRdy ),
       .io_deqRdy( T1603 ),
       .io_enqValid( T1602 ),
       .io_deqValid( fifo_42_io_deqValid ),
       .io_rst( T1601 )
  );
  fifo_0 fifo_43(.clk(clk), .reset(reset),
       .io_enqData( T1600 ),
       .io_deqData( fifo_43_io_deqData ),
       .io_enqRdy( fifo_43_io_enqRdy ),
       .io_deqRdy( T1599 ),
       .io_enqValid( T1598 ),
       .io_deqValid( fifo_43_io_deqValid ),
       .io_rst( T1597 )
  );
  fifo_0 fifo_44(.clk(clk), .reset(reset),
       .io_enqData( T1596 ),
       .io_deqData( fifo_44_io_deqData ),
       .io_enqRdy( fifo_44_io_enqRdy ),
       .io_deqRdy( T1595 ),
       .io_enqValid( T1594 ),
       .io_deqValid( fifo_44_io_deqValid ),
       .io_rst( T1593 )
  );
  fifo_0 fifo_45(.clk(clk), .reset(reset),
       .io_enqData( T1592 ),
       .io_deqData( fifo_45_io_deqData ),
       .io_enqRdy( fifo_45_io_enqRdy ),
       .io_deqRdy( T1591 ),
       .io_enqValid( T1590 ),
       .io_deqValid( fifo_45_io_deqValid ),
       .io_rst( T1589 )
  );
  fifo_0 fifo_46(.clk(clk), .reset(reset),
       .io_enqData( T1588 ),
       .io_deqData( fifo_46_io_deqData ),
       .io_enqRdy( fifo_46_io_enqRdy ),
       .io_deqRdy( T1587 ),
       .io_enqValid( T1586 ),
       .io_deqValid( fifo_46_io_deqValid ),
       .io_rst( T1585 )
  );
  fifo_0 fifo_47(.clk(clk), .reset(reset),
       .io_enqData( T1569 ),
       .io_deqData( fifo_47_io_deqData ),
       .io_enqRdy( fifo_47_io_enqRdy ),
       .io_deqRdy( T268 ),
       .io_enqValid( T1 ),
       .io_deqValid( fifo_47_io_deqValid ),
       .io_rst( T0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      nextSeqSelReg <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      nextSeqSelReg <= 1'h0;
    end else if(allDone) begin
      nextSeqSelReg <= T62;
    end
    if(reset) begin
      nextSeqReg2 <= 89'h0;
    end else if(T174) begin
      nextSeqReg2 <= nextSeqWire;
    end
    if(reset) begin
      firstSeqSelReg <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      firstSeqSelReg <= 1'h0;
    end else if(T177) begin
      firstSeqSelReg <= 1'h1;
    end
    if(reset) begin
      bankReadDoneReg_1 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_1 <= 1'h0;
    end else begin
      bankReadDoneReg_1 <= readDone_1;
    end
    if(reset) begin
      nextSeqRegValid2 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      nextSeqRegValid2 <= 1'h0;
    end else if(T195) begin
      nextSeqRegValid2 <= 1'h0;
    end else if(T194) begin
      nextSeqRegValid2 <= 1'h0;
    end else if(T174) begin
      nextSeqRegValid2 <= 1'h1;
    end
    if(reset) begin
      nextSeqRegValid1 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      nextSeqRegValid1 <= 1'h0;
    end else if(T177) begin
      nextSeqRegValid1 <= 1'h1;
    end
    if(reset) begin
      bankReadDoneReg_2 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_2 <= 1'h0;
    end else begin
      bankReadDoneReg_2 <= readDone_2;
    end
    if(reset) begin
      bankReadDoneReg_3 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_3 <= 1'h0;
    end else begin
      bankReadDoneReg_3 <= readDone_3;
    end
    if(reset) begin
      bankReadDoneReg_4 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_4 <= 1'h0;
    end else begin
      bankReadDoneReg_4 <= readDone_4;
    end
    if(reset) begin
      bankReadDoneReg_5 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_5 <= 1'h0;
    end else begin
      bankReadDoneReg_5 <= readDone_5;
    end
    if(reset) begin
      bankReadDoneReg_6 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_6 <= 1'h0;
    end else begin
      bankReadDoneReg_6 <= readDone_6;
    end
    if(reset) begin
      bankReadDoneReg_7 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_7 <= 1'h0;
    end else begin
      bankReadDoneReg_7 <= readDone_7;
    end
    if(reset) begin
      bankReadDoneReg_0 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      bankReadDoneReg_0 <= 1'h0;
    end else begin
      bankReadDoneReg_0 <= readDone_0;
    end
    if(reset) begin
      seqLevelDoneReg2 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      seqLevelDoneReg2 <= 1'h0;
    end else if(T1509) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1453) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1397) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1341) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1285) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1229) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1173) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1117) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1061) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T1005) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T949) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T893) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T837) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T781) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T725) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T669) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T613) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T557) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T501) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end else if(T361) begin
      seqLevelDoneReg2 <= seqLevelDoneReg1;
    end
    if(reset) begin
      bankSeqReg_0 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_1 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_2 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_3 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_4 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_5 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_6 <= 88'h0;
    end
    if(reset) begin
      bankSeqReg_7 <= 88'h0;
    end
    if(reset) begin
      seqLevelDoneReg1 <= 1'h0;
    end else if(fabInSeqMemConfig_io_rst) begin
      seqLevelDoneReg1 <= 1'h0;
    end else if(T67) begin
      seqLevelDoneReg1 <= T359;
    end else if(T78) begin
      seqLevelDoneReg1 <= T357;
    end else if(T89) begin
      seqLevelDoneReg1 <= T355;
    end else if(T100) begin
      seqLevelDoneReg1 <= T353;
    end else if(T111) begin
      seqLevelDoneReg1 <= T351;
    end else if(T122) begin
      seqLevelDoneReg1 <= T349;
    end else if(T133) begin
      seqLevelDoneReg1 <= T347;
    end else if(T143) begin
      seqLevelDoneReg1 <= T345;
    end
  end
endmodule

module fabInSeq(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_fabInData_19,
    output[31:0] io_fabInData_18,
    output[31:0] io_fabInData_17,
    output[31:0] io_fabInData_16,
    output[31:0] io_fabInData_15,
    output[31:0] io_fabInData_14,
    output[31:0] io_fabInData_13,
    output[31:0] io_fabInData_12,
    output[31:0] io_fabInData_11,
    output[31:0] io_fabInData_10,
    output[31:0] io_fabInData_9,
    output[31:0] io_fabInData_8,
    output[31:0] io_fabInData_7,
    output[31:0] io_fabInData_6,
    output[31:0] io_fabInData_5,
    output[31:0] io_fabInData_4,
    output[31:0] io_fabInData_3,
    output[31:0] io_fabInData_2,
    output[31:0] io_fabInData_1,
    output[31:0] io_fabInData_0,
    output io_fabInValid_19,
    output io_fabInValid_18,
    output io_fabInValid_17,
    output io_fabInValid_16,
    output io_fabInValid_15,
    output io_fabInValid_14,
    output io_fabInValid_13,
    output io_fabInValid_12,
    output io_fabInValid_11,
    output io_fabInValid_10,
    output io_fabInValid_9,
    output io_fabInValid_8,
    output io_fabInValid_7,
    output io_fabInValid_6,
    output io_fabInValid_5,
    output io_fabInValid_4,
    output io_fabInValid_3,
    output io_fabInValid_2,
    output io_fabInValid_1,
    output io_fabInValid_0,
    input  io_fabInRdy_19,
    input  io_fabInRdy_18,
    input  io_fabInRdy_17,
    input  io_fabInRdy_16,
    input  io_fabInRdy_15,
    input  io_fabInRdy_14,
    input  io_fabInRdy_13,
    input  io_fabInRdy_12,
    input  io_fabInRdy_11,
    input  io_fabInRdy_10,
    input  io_fabInRdy_9,
    input  io_fabInRdy_8,
    input  io_fabInRdy_7,
    input  io_fabInRdy_6,
    input  io_fabInRdy_5,
    input  io_fabInRdy_4,
    input  io_fabInRdy_3,
    input  io_fabInRdy_2,
    input  io_fabInRdy_1,
    input  io_fabInRdy_0,
    input [37:0] io_loadStore_7,
    input [37:0] io_loadStore_6,
    input [37:0] io_loadStore_5,
    input [37:0] io_loadStore_4,
    input [37:0] io_loadStore_3,
    input [37:0] io_loadStore_2,
    input [37:0] io_loadStore_1,
    input [37:0] io_loadStore_0,
    input  io_loadStoreValid_7,
    input  io_loadStoreValid_6,
    input  io_loadStoreValid_5,
    input  io_loadStoreValid_4,
    input  io_loadStoreValid_3,
    input  io_loadStoreValid_2,
    input  io_loadStoreValid_1,
    input  io_loadStoreValid_0,
    output io_loadStoreRdy_7,
    output io_loadStoreRdy_6,
    output io_loadStoreRdy_5,
    output io_loadStoreRdy_4,
    output io_loadStoreRdy_3,
    output io_loadStoreRdy_2,
    output io_loadStoreRdy_1,
    output io_loadStoreRdy_0,
    input [37:0] io_fabStore_7,
    input [37:0] io_fabStore_6,
    input [37:0] io_fabStore_5,
    input [37:0] io_fabStore_4,
    input [37:0] io_fabStore_3,
    input [37:0] io_fabStore_2,
    input [37:0] io_fabStore_1,
    input [37:0] io_fabStore_0,
    input  io_fabStoreValid_7,
    input  io_fabStoreValid_6,
    input  io_fabStoreValid_5,
    input  io_fabStoreValid_4,
    input  io_fabStoreValid_3,
    input  io_fabStoreValid_2,
    input  io_fabStoreValid_1,
    input  io_fabStoreValid_0,
    output io_fabStoreRdy_7,
    output io_fabStoreRdy_6,
    output io_fabStoreRdy_5,
    output io_fabStoreRdy_4,
    output io_fabStoreRdy_3,
    output io_fabStoreRdy_2,
    output io_fabStoreRdy_1,
    output io_fabStoreRdy_0,
    output io_computeDone
);

  wire[8:0] ctrlClass_io_seqMemAddr;
  wire ctrlClass_io_seqMemAddrValid;
  wire ctrlClass_io_computeDone;
  wire[31:0] dpClass_io_fabInData_19;
  wire[31:0] dpClass_io_fabInData_18;
  wire[31:0] dpClass_io_fabInData_17;
  wire[31:0] dpClass_io_fabInData_16;
  wire[31:0] dpClass_io_fabInData_15;
  wire[31:0] dpClass_io_fabInData_14;
  wire[31:0] dpClass_io_fabInData_13;
  wire[31:0] dpClass_io_fabInData_12;
  wire[31:0] dpClass_io_fabInData_11;
  wire[31:0] dpClass_io_fabInData_10;
  wire[31:0] dpClass_io_fabInData_9;
  wire[31:0] dpClass_io_fabInData_8;
  wire[31:0] dpClass_io_fabInData_7;
  wire[31:0] dpClass_io_fabInData_6;
  wire[31:0] dpClass_io_fabInData_5;
  wire[31:0] dpClass_io_fabInData_4;
  wire[31:0] dpClass_io_fabInData_3;
  wire[31:0] dpClass_io_fabInData_2;
  wire[31:0] dpClass_io_fabInData_1;
  wire[31:0] dpClass_io_fabInData_0;
  wire dpClass_io_fabInValid_19;
  wire dpClass_io_fabInValid_18;
  wire dpClass_io_fabInValid_17;
  wire dpClass_io_fabInValid_16;
  wire dpClass_io_fabInValid_15;
  wire dpClass_io_fabInValid_14;
  wire dpClass_io_fabInValid_13;
  wire dpClass_io_fabInValid_12;
  wire dpClass_io_fabInValid_11;
  wire dpClass_io_fabInValid_10;
  wire dpClass_io_fabInValid_9;
  wire dpClass_io_fabInValid_8;
  wire dpClass_io_fabInValid_7;
  wire dpClass_io_fabInValid_6;
  wire dpClass_io_fabInValid_5;
  wire dpClass_io_fabInValid_4;
  wire dpClass_io_fabInValid_3;
  wire dpClass_io_fabInValid_2;
  wire dpClass_io_fabInValid_1;
  wire dpClass_io_fabInValid_0;
  wire dpClass_io_loadStoreRdy_7;
  wire dpClass_io_loadStoreRdy_6;
  wire dpClass_io_loadStoreRdy_5;
  wire dpClass_io_loadStoreRdy_4;
  wire dpClass_io_loadStoreRdy_3;
  wire dpClass_io_loadStoreRdy_2;
  wire dpClass_io_loadStoreRdy_1;
  wire dpClass_io_loadStoreRdy_0;
  wire dpClass_io_fabStoreRdy_7;
  wire dpClass_io_fabStoreRdy_6;
  wire dpClass_io_fabStoreRdy_5;
  wire dpClass_io_fabStoreRdy_4;
  wire dpClass_io_fabStoreRdy_3;
  wire dpClass_io_fabStoreRdy_2;
  wire dpClass_io_fabStoreRdy_1;
  wire dpClass_io_fabStoreRdy_0;
  wire dpClass_io_seqProceed;


  assign io_computeDone = ctrlClass_io_computeDone;
  assign io_fabStoreRdy_0 = dpClass_io_fabStoreRdy_0;
  assign io_fabStoreRdy_1 = dpClass_io_fabStoreRdy_1;
  assign io_fabStoreRdy_2 = dpClass_io_fabStoreRdy_2;
  assign io_fabStoreRdy_3 = dpClass_io_fabStoreRdy_3;
  assign io_fabStoreRdy_4 = dpClass_io_fabStoreRdy_4;
  assign io_fabStoreRdy_5 = dpClass_io_fabStoreRdy_5;
  assign io_fabStoreRdy_6 = dpClass_io_fabStoreRdy_6;
  assign io_fabStoreRdy_7 = dpClass_io_fabStoreRdy_7;
  assign io_loadStoreRdy_0 = dpClass_io_loadStoreRdy_0;
  assign io_loadStoreRdy_1 = dpClass_io_loadStoreRdy_1;
  assign io_loadStoreRdy_2 = dpClass_io_loadStoreRdy_2;
  assign io_loadStoreRdy_3 = dpClass_io_loadStoreRdy_3;
  assign io_loadStoreRdy_4 = dpClass_io_loadStoreRdy_4;
  assign io_loadStoreRdy_5 = dpClass_io_loadStoreRdy_5;
  assign io_loadStoreRdy_6 = dpClass_io_loadStoreRdy_6;
  assign io_loadStoreRdy_7 = dpClass_io_loadStoreRdy_7;
  assign io_fabInValid_0 = dpClass_io_fabInValid_0;
  assign io_fabInValid_1 = dpClass_io_fabInValid_1;
  assign io_fabInValid_2 = dpClass_io_fabInValid_2;
  assign io_fabInValid_3 = dpClass_io_fabInValid_3;
  assign io_fabInValid_4 = dpClass_io_fabInValid_4;
  assign io_fabInValid_5 = dpClass_io_fabInValid_5;
  assign io_fabInValid_6 = dpClass_io_fabInValid_6;
  assign io_fabInValid_7 = dpClass_io_fabInValid_7;
  assign io_fabInValid_8 = dpClass_io_fabInValid_8;
  assign io_fabInValid_9 = dpClass_io_fabInValid_9;
  assign io_fabInValid_10 = dpClass_io_fabInValid_10;
  assign io_fabInValid_11 = dpClass_io_fabInValid_11;
  assign io_fabInValid_12 = dpClass_io_fabInValid_12;
  assign io_fabInValid_13 = dpClass_io_fabInValid_13;
  assign io_fabInValid_14 = dpClass_io_fabInValid_14;
  assign io_fabInValid_15 = dpClass_io_fabInValid_15;
  assign io_fabInValid_16 = dpClass_io_fabInValid_16;
  assign io_fabInValid_17 = dpClass_io_fabInValid_17;
  assign io_fabInValid_18 = dpClass_io_fabInValid_18;
  assign io_fabInValid_19 = dpClass_io_fabInValid_19;
  assign io_fabInData_0 = dpClass_io_fabInData_0;
  assign io_fabInData_1 = dpClass_io_fabInData_1;
  assign io_fabInData_2 = dpClass_io_fabInData_2;
  assign io_fabInData_3 = dpClass_io_fabInData_3;
  assign io_fabInData_4 = dpClass_io_fabInData_4;
  assign io_fabInData_5 = dpClass_io_fabInData_5;
  assign io_fabInData_6 = dpClass_io_fabInData_6;
  assign io_fabInData_7 = dpClass_io_fabInData_7;
  assign io_fabInData_8 = dpClass_io_fabInData_8;
  assign io_fabInData_9 = dpClass_io_fabInData_9;
  assign io_fabInData_10 = dpClass_io_fabInData_10;
  assign io_fabInData_11 = dpClass_io_fabInData_11;
  assign io_fabInData_12 = dpClass_io_fabInData_12;
  assign io_fabInData_13 = dpClass_io_fabInData_13;
  assign io_fabInData_14 = dpClass_io_fabInData_14;
  assign io_fabInData_15 = dpClass_io_fabInData_15;
  assign io_fabInData_16 = dpClass_io_fabInData_16;
  assign io_fabInData_17 = dpClass_io_fabInData_17;
  assign io_fabInData_18 = dpClass_io_fabInData_18;
  assign io_fabInData_19 = dpClass_io_fabInData_19;
  fabInSeqCtrl ctrlClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( ctrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( ctrlClass_io_seqMemAddrValid ),
       .io_seqProceed( dpClass_io_seqProceed ),
       .io_computeDone( ctrlClass_io_computeDone )
  );
  fabInSeqDP dpClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( ctrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( ctrlClass_io_seqMemAddrValid ),
       .io_fabInData_19( dpClass_io_fabInData_19 ),
       .io_fabInData_18( dpClass_io_fabInData_18 ),
       .io_fabInData_17( dpClass_io_fabInData_17 ),
       .io_fabInData_16( dpClass_io_fabInData_16 ),
       .io_fabInData_15( dpClass_io_fabInData_15 ),
       .io_fabInData_14( dpClass_io_fabInData_14 ),
       .io_fabInData_13( dpClass_io_fabInData_13 ),
       .io_fabInData_12( dpClass_io_fabInData_12 ),
       .io_fabInData_11( dpClass_io_fabInData_11 ),
       .io_fabInData_10( dpClass_io_fabInData_10 ),
       .io_fabInData_9( dpClass_io_fabInData_9 ),
       .io_fabInData_8( dpClass_io_fabInData_8 ),
       .io_fabInData_7( dpClass_io_fabInData_7 ),
       .io_fabInData_6( dpClass_io_fabInData_6 ),
       .io_fabInData_5( dpClass_io_fabInData_5 ),
       .io_fabInData_4( dpClass_io_fabInData_4 ),
       .io_fabInData_3( dpClass_io_fabInData_3 ),
       .io_fabInData_2( dpClass_io_fabInData_2 ),
       .io_fabInData_1( dpClass_io_fabInData_1 ),
       .io_fabInData_0( dpClass_io_fabInData_0 ),
       .io_fabInValid_19( dpClass_io_fabInValid_19 ),
       .io_fabInValid_18( dpClass_io_fabInValid_18 ),
       .io_fabInValid_17( dpClass_io_fabInValid_17 ),
       .io_fabInValid_16( dpClass_io_fabInValid_16 ),
       .io_fabInValid_15( dpClass_io_fabInValid_15 ),
       .io_fabInValid_14( dpClass_io_fabInValid_14 ),
       .io_fabInValid_13( dpClass_io_fabInValid_13 ),
       .io_fabInValid_12( dpClass_io_fabInValid_12 ),
       .io_fabInValid_11( dpClass_io_fabInValid_11 ),
       .io_fabInValid_10( dpClass_io_fabInValid_10 ),
       .io_fabInValid_9( dpClass_io_fabInValid_9 ),
       .io_fabInValid_8( dpClass_io_fabInValid_8 ),
       .io_fabInValid_7( dpClass_io_fabInValid_7 ),
       .io_fabInValid_6( dpClass_io_fabInValid_6 ),
       .io_fabInValid_5( dpClass_io_fabInValid_5 ),
       .io_fabInValid_4( dpClass_io_fabInValid_4 ),
       .io_fabInValid_3( dpClass_io_fabInValid_3 ),
       .io_fabInValid_2( dpClass_io_fabInValid_2 ),
       .io_fabInValid_1( dpClass_io_fabInValid_1 ),
       .io_fabInValid_0( dpClass_io_fabInValid_0 ),
       .io_fabInRdy_19( io_fabInRdy_19 ),
       .io_fabInRdy_18( io_fabInRdy_18 ),
       .io_fabInRdy_17( io_fabInRdy_17 ),
       .io_fabInRdy_16( io_fabInRdy_16 ),
       .io_fabInRdy_15( io_fabInRdy_15 ),
       .io_fabInRdy_14( io_fabInRdy_14 ),
       .io_fabInRdy_13( io_fabInRdy_13 ),
       .io_fabInRdy_12( io_fabInRdy_12 ),
       .io_fabInRdy_11( io_fabInRdy_11 ),
       .io_fabInRdy_10( io_fabInRdy_10 ),
       .io_fabInRdy_9( io_fabInRdy_9 ),
       .io_fabInRdy_8( io_fabInRdy_8 ),
       .io_fabInRdy_7( io_fabInRdy_7 ),
       .io_fabInRdy_6( io_fabInRdy_6 ),
       .io_fabInRdy_5( io_fabInRdy_5 ),
       .io_fabInRdy_4( io_fabInRdy_4 ),
       .io_fabInRdy_3( io_fabInRdy_3 ),
       .io_fabInRdy_2( io_fabInRdy_2 ),
       .io_fabInRdy_1( io_fabInRdy_1 ),
       .io_fabInRdy_0( io_fabInRdy_0 ),
       .io_loadStore_7( io_loadStore_7 ),
       .io_loadStore_6( io_loadStore_6 ),
       .io_loadStore_5( io_loadStore_5 ),
       .io_loadStore_4( io_loadStore_4 ),
       .io_loadStore_3( io_loadStore_3 ),
       .io_loadStore_2( io_loadStore_2 ),
       .io_loadStore_1( io_loadStore_1 ),
       .io_loadStore_0( io_loadStore_0 ),
       .io_loadStoreValid_7( io_loadStoreValid_7 ),
       .io_loadStoreValid_6( io_loadStoreValid_6 ),
       .io_loadStoreValid_5( io_loadStoreValid_5 ),
       .io_loadStoreValid_4( io_loadStoreValid_4 ),
       .io_loadStoreValid_3( io_loadStoreValid_3 ),
       .io_loadStoreValid_2( io_loadStoreValid_2 ),
       .io_loadStoreValid_1( io_loadStoreValid_1 ),
       .io_loadStoreValid_0( io_loadStoreValid_0 ),
       .io_loadStoreRdy_7( dpClass_io_loadStoreRdy_7 ),
       .io_loadStoreRdy_6( dpClass_io_loadStoreRdy_6 ),
       .io_loadStoreRdy_5( dpClass_io_loadStoreRdy_5 ),
       .io_loadStoreRdy_4( dpClass_io_loadStoreRdy_4 ),
       .io_loadStoreRdy_3( dpClass_io_loadStoreRdy_3 ),
       .io_loadStoreRdy_2( dpClass_io_loadStoreRdy_2 ),
       .io_loadStoreRdy_1( dpClass_io_loadStoreRdy_1 ),
       .io_loadStoreRdy_0( dpClass_io_loadStoreRdy_0 ),
       .io_fabStore_7( io_fabStore_7 ),
       .io_fabStore_6( io_fabStore_6 ),
       .io_fabStore_5( io_fabStore_5 ),
       .io_fabStore_4( io_fabStore_4 ),
       .io_fabStore_3( io_fabStore_3 ),
       .io_fabStore_2( io_fabStore_2 ),
       .io_fabStore_1( io_fabStore_1 ),
       .io_fabStore_0( io_fabStore_0 ),
       .io_fabStoreValid_7( io_fabStoreValid_7 ),
       .io_fabStoreValid_6( io_fabStoreValid_6 ),
       .io_fabStoreValid_5( io_fabStoreValid_5 ),
       .io_fabStoreValid_4( io_fabStoreValid_4 ),
       .io_fabStoreValid_3( io_fabStoreValid_3 ),
       .io_fabStoreValid_2( io_fabStoreValid_2 ),
       .io_fabStoreValid_1( io_fabStoreValid_1 ),
       .io_fabStoreValid_0( io_fabStoreValid_0 ),
       .io_fabStoreRdy_7( dpClass_io_fabStoreRdy_7 ),
       .io_fabStoreRdy_6( dpClass_io_fabStoreRdy_6 ),
       .io_fabStoreRdy_5( dpClass_io_fabStoreRdy_5 ),
       .io_fabStoreRdy_4( dpClass_io_fabStoreRdy_4 ),
       .io_fabStoreRdy_3( dpClass_io_fabStoreRdy_3 ),
       .io_fabStoreRdy_2( dpClass_io_fabStoreRdy_2 ),
       .io_fabStoreRdy_1( dpClass_io_fabStoreRdy_1 ),
       .io_fabStoreRdy_0( dpClass_io_fabStoreRdy_0 ),
       .io_seqProceed( dpClass_io_seqProceed )
  );
endmodule

module fabOutSeqCtrl(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input  io_outLocValid_19,
    input  io_outLocValid_18,
    input  io_outLocValid_17,
    input  io_outLocValid_16,
    input  io_outLocValid_15,
    input  io_outLocValid_14,
    input  io_outLocValid_13,
    input  io_outLocValid_12,
    input  io_outLocValid_11,
    input  io_outLocValid_10,
    input  io_outLocValid_9,
    input  io_outLocValid_8,
    input  io_outLocValid_7,
    input  io_outLocValid_6,
    input  io_outLocValid_5,
    input  io_outLocValid_4,
    input  io_outLocValid_3,
    input  io_outLocValid_2,
    input  io_outLocValid_1,
    input  io_outLocValid_0,
    output[8:0] io_seqMemAddr_19,
    output[8:0] io_seqMemAddr_18,
    output[8:0] io_seqMemAddr_17,
    output[8:0] io_seqMemAddr_16,
    output[8:0] io_seqMemAddr_15,
    output[8:0] io_seqMemAddr_14,
    output[8:0] io_seqMemAddr_13,
    output[8:0] io_seqMemAddr_12,
    output[8:0] io_seqMemAddr_11,
    output[8:0] io_seqMemAddr_10,
    output[8:0] io_seqMemAddr_9,
    output[8:0] io_seqMemAddr_8,
    output[8:0] io_seqMemAddr_7,
    output[8:0] io_seqMemAddr_6,
    output[8:0] io_seqMemAddr_5,
    output[8:0] io_seqMemAddr_4,
    output[8:0] io_seqMemAddr_3,
    output[8:0] io_seqMemAddr_2,
    output[8:0] io_seqMemAddr_1,
    output[8:0] io_seqMemAddr_0,
    output io_seqMemAddrValid_19,
    output io_seqMemAddrValid_18,
    output io_seqMemAddrValid_17,
    output io_seqMemAddrValid_16,
    output io_seqMemAddrValid_15,
    output io_seqMemAddrValid_14,
    output io_seqMemAddrValid_13,
    output io_seqMemAddrValid_12,
    output io_seqMemAddrValid_11,
    output io_seqMemAddrValid_10,
    output io_seqMemAddrValid_9,
    output io_seqMemAddrValid_8,
    output io_seqMemAddrValid_7,
    output io_seqMemAddrValid_6,
    output io_seqMemAddrValid_5,
    output io_seqMemAddrValid_4,
    output io_seqMemAddrValid_3,
    output io_seqMemAddrValid_2,
    output io_seqMemAddrValid_1,
    output io_seqMemAddrValid_0,
    input  io_seqProceed_19,
    input  io_seqProceed_18,
    input  io_seqProceed_17,
    input  io_seqProceed_16,
    input  io_seqProceed_15,
    input  io_seqProceed_14,
    input  io_seqProceed_13,
    input  io_seqProceed_12,
    input  io_seqProceed_11,
    input  io_seqProceed_10,
    input  io_seqProceed_9,
    input  io_seqProceed_8,
    input  io_seqProceed_7,
    input  io_seqProceed_6,
    input  io_seqProceed_5,
    input  io_seqProceed_4,
    input  io_seqProceed_3,
    input  io_seqProceed_2,
    input  io_seqProceed_1,
    input  io_seqProceed_0
);

  wire T0;
  wire T1;
  reg  computeEnable;
  wire T1645;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[514:0] lastAddr;
  wire[514:0] T1646;
  wire[513:0] T8;
  wire[513:0] T1647;
  reg [8:0] epilogueDepth;
  wire[8:0] T1648;
  wire[8:0] T9;
  wire[8:0] T1649;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire[9:0] T23;
  wire[513:0] ssEnd;
  wire[513:0] T1650;
  wire[8:0] T24;
  reg [8:0] steadyStateDepth;
  wire[8:0] T1651;
  wire[9:0] T1652;
  wire[9:0] T25;
  wire[9:0] T1653;
  wire[9:0] T26;
  wire T27;
  reg [8:0] prologueDepth;
  wire[8:0] T1654;
  wire[8:0] T28;
  wire[8:0] T1655;
  wire[6:0] T29;
  wire startComputeValid;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire computeDone;
  wire T34;
  wire T35;
  wire resetComputeValid;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg  reqDone_0;
  wire T1656;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire reqDoneWire_19;
  wire T88;
  wire T89;
  wire T90;
  wire T131;
  wire T132;
  wire T133;
  wire nextRequest_19;
  wire T134;
  wire T135;
  reg  reqDone_19;
  wire T1657;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T136;
  wire T137;
  wire T138;
  wire reqDoneWire_18;
  wire T139;
  wire T140;
  wire T141;
  wire T182;
  wire T183;
  wire T184;
  wire nextRequest_18;
  wire T185;
  wire T186;
  reg  reqDone_18;
  wire T1658;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T187;
  wire T188;
  wire T189;
  wire reqDoneWire_17;
  wire T190;
  wire T191;
  wire T192;
  wire T233;
  wire T234;
  wire T235;
  wire nextRequest_17;
  wire T236;
  wire T237;
  reg  reqDone_17;
  wire T1659;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T238;
  wire T239;
  wire T240;
  wire reqDoneWire_16;
  wire T241;
  wire T242;
  wire T243;
  wire T284;
  wire T285;
  wire T286;
  wire nextRequest_16;
  wire T287;
  wire T288;
  reg  reqDone_16;
  wire T1660;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T289;
  wire T290;
  wire T291;
  wire reqDoneWire_15;
  wire T292;
  wire T293;
  wire T294;
  wire T335;
  wire T336;
  wire T337;
  wire nextRequest_15;
  wire T338;
  wire T339;
  reg  reqDone_15;
  wire T1661;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T340;
  wire T341;
  wire T342;
  wire reqDoneWire_14;
  wire T343;
  wire T344;
  wire T345;
  wire T386;
  wire T387;
  wire T388;
  wire nextRequest_14;
  wire T389;
  wire T390;
  reg  reqDone_14;
  wire T1662;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T391;
  wire T392;
  wire T393;
  wire reqDoneWire_13;
  wire T394;
  wire T395;
  wire T396;
  wire T437;
  wire T438;
  wire T439;
  wire nextRequest_13;
  wire T440;
  wire T441;
  reg  reqDone_13;
  wire T1663;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T442;
  wire T443;
  wire T444;
  wire reqDoneWire_12;
  wire T445;
  wire T446;
  wire T447;
  wire T488;
  wire T489;
  wire T490;
  wire nextRequest_12;
  wire T491;
  wire T492;
  reg  reqDone_12;
  wire T1664;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T493;
  wire T494;
  wire T495;
  wire reqDoneWire_11;
  wire T496;
  wire T497;
  wire T498;
  wire T539;
  wire T540;
  wire T541;
  wire nextRequest_11;
  wire T542;
  wire T543;
  reg  reqDone_11;
  wire T1665;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T544;
  wire T545;
  wire T546;
  wire reqDoneWire_10;
  wire T547;
  wire T548;
  wire T549;
  wire T590;
  wire T591;
  wire T592;
  wire nextRequest_10;
  wire T593;
  wire T594;
  reg  reqDone_10;
  wire T1666;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T595;
  wire T596;
  wire T597;
  wire reqDoneWire_9;
  wire T598;
  wire T599;
  wire T600;
  wire T641;
  wire T642;
  wire T643;
  wire nextRequest_9;
  wire T644;
  wire T645;
  reg  reqDone_9;
  wire T1667;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T646;
  wire T647;
  wire T648;
  wire reqDoneWire_8;
  wire T649;
  wire T650;
  wire T651;
  wire T692;
  wire T693;
  wire T694;
  wire nextRequest_8;
  wire T695;
  wire T696;
  reg  reqDone_8;
  wire T1668;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T697;
  wire T698;
  wire T699;
  wire reqDoneWire_7;
  wire T700;
  wire T701;
  wire T702;
  wire T743;
  wire T744;
  wire T745;
  wire nextRequest_7;
  wire T746;
  wire T747;
  reg  reqDone_7;
  wire T1669;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T748;
  wire T749;
  wire T750;
  wire reqDoneWire_6;
  wire T751;
  wire T752;
  wire T753;
  wire T794;
  wire T795;
  wire T796;
  wire nextRequest_6;
  wire T797;
  wire T798;
  reg  reqDone_6;
  wire T1670;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T799;
  wire T800;
  wire T801;
  wire reqDoneWire_5;
  wire T802;
  wire T803;
  wire T804;
  wire T845;
  wire T846;
  wire T847;
  wire nextRequest_5;
  wire T848;
  wire T849;
  reg  reqDone_5;
  wire T1671;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T850;
  wire T851;
  wire T852;
  wire reqDoneWire_4;
  wire T853;
  wire T854;
  wire T855;
  wire T896;
  wire T897;
  wire T898;
  wire nextRequest_4;
  wire T899;
  wire T900;
  reg  reqDone_4;
  wire T1672;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T901;
  wire T902;
  wire T903;
  wire reqDoneWire_3;
  wire T904;
  wire T905;
  wire T906;
  wire T947;
  wire T948;
  wire T949;
  wire nextRequest_3;
  wire T950;
  wire T951;
  reg  reqDone_3;
  wire T1673;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T952;
  wire T953;
  wire T954;
  wire reqDoneWire_2;
  wire T955;
  wire T956;
  wire T957;
  wire T998;
  wire T999;
  wire T1000;
  wire nextRequest_2;
  wire T1001;
  wire T1002;
  reg  reqDone_2;
  wire T1674;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T1003;
  wire T1004;
  wire T1005;
  wire reqDoneWire_1;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1049;
  wire T1050;
  wire T1051;
  wire nextRequest_1;
  wire T1052;
  wire T1053;
  reg  reqDone_1;
  wire T1675;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1054;
  wire T1055;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire reqDoneWire_0;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire nextRequest_0;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1484;
  wire T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire T1497;
  wire T1498;
  wire T1499;
  wire T1500;
  wire T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire T1508;
  wire T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire T1516;
  wire T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire T1540;
  wire T1541;
  wire T1542;
  wire[8:0] T1543;
  reg [8:0] seqMemAddr;
  wire[8:0] T1676;
  wire[513:0] T1677;
  wire[513:0] T1544;
  wire[513:0] T1545;
  wire[513:0] T1678;
  wire[8:0] T1546;
  wire[8:0] T1547;
  wire[8:0] T1548;
  wire T1549;
  wire T1550;
  wire nextSeqRdy;
  wire T1551;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire T1556;
  wire T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire T1577;
  wire T1578;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire T1585;
  wire T1586;
  wire T1587;
  wire T1588;
  wire T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  reg [8:0] epilogueSpill;
  wire[8:0] T1679;
  wire[9:0] T1680;
  wire[9:0] T1593;
  wire[9:0] T1681;
  wire[9:0] T1594;
  wire T1595;
  wire[31:0] T1596;
  reg [31:0] iterCount;
  wire[31:0] T1682;
  wire[31:0] T1597;
  wire[31:0] T1683;
  wire[18:0] T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire[2:0] T1602;
  wire T1603;
  reg [31:0] currentIter;
  wire[31:0] T1684;
  wire[31:0] T1604;
  wire[31:0] T1605;
  wire[31:0] T1606;
  wire T1607;
  wire T1608;
  wire[513:0] T1609;
  wire[513:0] T1685;
  wire T1610;
  wire T1611;
  wire[8:0] T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire[513:0] T1619;
  wire[513:0] T1686;
  wire T1620;
  wire T1621;
  wire[513:0] T1687;
  wire[8:0] T1622;
  wire T1623;
  wire T1624;
  wire T1625;
  wire[8:0] T1626;
  wire[8:0] T1627;
  wire[8:0] T1628;
  wire[8:0] T1629;
  wire[8:0] T1630;
  wire[8:0] T1631;
  wire[8:0] T1632;
  wire[8:0] T1633;
  wire[8:0] T1634;
  wire[8:0] T1635;
  wire[8:0] T1636;
  wire[8:0] T1637;
  wire[8:0] T1638;
  wire[8:0] T1639;
  wire[8:0] T1640;
  wire[8:0] T1641;
  wire[8:0] T1642;
  wire[8:0] T1643;
  wire[8:0] T1644;
  wire fabOutSeqCtrlConfigure_io_computeCtrl;
  wire fabOutSeqCtrlConfigure_io_computeCtrlValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    computeEnable = {1{$random}};
    epilogueDepth = {1{$random}};
    steadyStateDepth = {1{$random}};
    prologueDepth = {1{$random}};
    reqDone_0 = {1{$random}};
    reqDone_19 = {1{$random}};
    reqDone_18 = {1{$random}};
    reqDone_17 = {1{$random}};
    reqDone_16 = {1{$random}};
    reqDone_15 = {1{$random}};
    reqDone_14 = {1{$random}};
    reqDone_13 = {1{$random}};
    reqDone_12 = {1{$random}};
    reqDone_11 = {1{$random}};
    reqDone_10 = {1{$random}};
    reqDone_9 = {1{$random}};
    reqDone_8 = {1{$random}};
    reqDone_7 = {1{$random}};
    reqDone_6 = {1{$random}};
    reqDone_5 = {1{$random}};
    reqDone_4 = {1{$random}};
    reqDone_3 = {1{$random}};
    reqDone_2 = {1{$random}};
    reqDone_1 = {1{$random}};
    seqMemAddr = {1{$random}};
    epilogueSpill = {1{$random}};
    iterCount = {1{$random}};
    currentIter = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_seqMemAddrValid_0 = T0;
  assign T0 = T1 ? 1'h1 : 1'h0;
  assign T1 = T45 & computeEnable;
  assign T1645 = reset ? 1'h0 : T2;
  assign T2 = T42 ? 1'h0 : T3;
  assign T3 = T39 ? 1'h0 : T4;
  assign T4 = T5 ? 1'h1 : computeEnable;
  assign T5 = T33 & T6;
  assign T6 = startComputeValid & T7;
  assign T7 = lastAddr != 515'h0;
  assign lastAddr = T1646;
  assign T1646 = {1'h0, T8};
  assign T8 = ssEnd + T1647;
  assign T1647 = {505'h0, epilogueDepth};
  assign T1648 = reset ? 9'h0 : T9;
  assign T9 = T11 ? T1649 : epilogueDepth;
  assign T1649 = {2'h0, T10};
  assign T10 = io_inConfig[3'h6:1'h0];
  assign T11 = T18 & T12;
  assign T12 = T15 & T13;
  assign T13 = T14 == 1'h1;
  assign T14 = io_inConfig[5'h11:5'h11];
  assign T15 = T16 ^ 1'h1;
  assign T16 = T17 == 1'h0;
  assign T17 = io_inConfig[5'h11:5'h11];
  assign T18 = T21 & T19;
  assign T19 = T20 == 3'h0;
  assign T20 = io_inConfig[5'h15:5'h13];
  assign T21 = io_inValid & T22;
  assign T22 = T23 == 10'h102;
  assign T23 = io_inConfig[5'h1f:5'h16];
  assign ssEnd = T1650;
  assign T1650 = {505'h0, T24};
  assign T24 = prologueDepth + steadyStateDepth;
  assign T1651 = T1652[4'h8:1'h0];
  assign T1652 = reset ? 10'h0 : T25;
  assign T25 = T27 ? T26 : T1653;
  assign T1653 = {1'h0, steadyStateDepth};
  assign T26 = io_inConfig[5'h10:3'h7];
  assign T27 = T18 & T16;
  assign T1654 = reset ? 9'h0 : T28;
  assign T28 = T27 ? T1655 : prologueDepth;
  assign T1655 = {2'h0, T29};
  assign T29 = io_inConfig[3'h6:1'h0];
  assign startComputeValid = T30;
  assign T30 = T32 ? 1'h0 : T31;
  assign T31 = fabOutSeqCtrlConfigure_io_computeCtrlValid & fabOutSeqCtrlConfigure_io_computeCtrl;
  assign T32 = fabOutSeqCtrlConfigure_io_computeCtrlValid ^ 1'h1;
  assign T33 = T35 | computeDone;
  assign computeDone = T34;
  assign T34 = computeEnable ^ 1'h1;
  assign T35 = startComputeValid | resetComputeValid;
  assign resetComputeValid = T36;
  assign T36 = T32 ? 1'h0 : T37;
  assign T37 = fabOutSeqCtrlConfigure_io_computeCtrlValid & T38;
  assign T38 = fabOutSeqCtrlConfigure_io_computeCtrl ^ 1'h1;
  assign T39 = T33 & T40;
  assign T40 = T41 & resetComputeValid;
  assign T41 = T6 ^ 1'h1;
  assign T42 = T33 & T43;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T6 | resetComputeValid;
  assign T45 = ~ reqDone_0;
  assign T1656 = reset ? 1'h0 : T46;
  assign T46 = T1484 ? reqDoneWire_0 : T47;
  assign T47 = T1464 ? 1'h0 : T48;
  assign T48 = T1462 ? reqDoneWire_0 : T49;
  assign T49 = T1442 ? 1'h0 : T50;
  assign T50 = T1440 ? reqDoneWire_0 : T51;
  assign T51 = T1420 ? 1'h0 : T52;
  assign T52 = T1418 ? reqDoneWire_0 : T53;
  assign T53 = T1398 ? 1'h0 : T54;
  assign T54 = T1396 ? reqDoneWire_0 : T55;
  assign T55 = T1376 ? 1'h0 : T56;
  assign T56 = T1374 ? reqDoneWire_0 : T57;
  assign T57 = T1354 ? 1'h0 : T58;
  assign T58 = T1352 ? reqDoneWire_0 : T59;
  assign T59 = T1332 ? 1'h0 : T60;
  assign T60 = T1330 ? reqDoneWire_0 : T61;
  assign T61 = T1310 ? 1'h0 : T62;
  assign T62 = T1308 ? reqDoneWire_0 : T63;
  assign T63 = T1288 ? 1'h0 : T64;
  assign T64 = T1286 ? reqDoneWire_0 : T65;
  assign T65 = T1266 ? 1'h0 : T66;
  assign T66 = T1264 ? reqDoneWire_0 : T67;
  assign T67 = T1244 ? 1'h0 : T68;
  assign T68 = T1242 ? reqDoneWire_0 : T69;
  assign T69 = T1222 ? 1'h0 : T70;
  assign T70 = T1220 ? reqDoneWire_0 : T71;
  assign T71 = T1200 ? 1'h0 : T72;
  assign T72 = T1198 ? reqDoneWire_0 : T73;
  assign T73 = T1178 ? 1'h0 : T74;
  assign T74 = T1176 ? reqDoneWire_0 : T75;
  assign T75 = T1156 ? 1'h0 : T76;
  assign T76 = T1154 ? reqDoneWire_0 : T77;
  assign T77 = T1134 ? 1'h0 : T78;
  assign T78 = T1132 ? reqDoneWire_0 : T79;
  assign T79 = T1112 ? 1'h0 : T80;
  assign T80 = T1110 ? reqDoneWire_0 : T81;
  assign T81 = T1090 ? 1'h0 : T82;
  assign T82 = T1088 ? reqDoneWire_0 : T83;
  assign T83 = T1068 ? 1'h0 : T84;
  assign T84 = T1066 ? reqDoneWire_0 : T85;
  assign T85 = T86 ? 1'h0 : reqDone_0;
  assign T86 = computeEnable & T87;
  assign T87 = T138 & reqDoneWire_19;
  assign reqDoneWire_19 = T88;
  assign T88 = T136 ? reqDone_19 : T89;
  assign T89 = T131 ? 1'h1 : T90;
  assign T90 = computeEnable ? reqDone_19 : 1'h0;
  assign T131 = computeEnable & T132;
  assign T132 = nextRequest_19 | T133;
  assign T133 = ~ io_outLocValid_19;
  assign nextRequest_19 = T134;
  assign T134 = T135 ? 1'h0 : io_seqProceed_19;
  assign T135 = io_seqProceed_19 ^ 1'h1;
  assign T1657 = reset ? 1'h0 : T91;
  assign T91 = T1484 ? reqDoneWire_19 : T92;
  assign T92 = T1464 ? 1'h0 : T93;
  assign T93 = T1462 ? reqDoneWire_19 : T94;
  assign T94 = T1442 ? 1'h0 : T95;
  assign T95 = T1440 ? reqDoneWire_19 : T96;
  assign T96 = T1420 ? 1'h0 : T97;
  assign T97 = T1418 ? reqDoneWire_19 : T98;
  assign T98 = T1398 ? 1'h0 : T99;
  assign T99 = T1396 ? reqDoneWire_19 : T100;
  assign T100 = T1376 ? 1'h0 : T101;
  assign T101 = T1374 ? reqDoneWire_19 : T102;
  assign T102 = T1354 ? 1'h0 : T103;
  assign T103 = T1352 ? reqDoneWire_19 : T104;
  assign T104 = T1332 ? 1'h0 : T105;
  assign T105 = T1330 ? reqDoneWire_19 : T106;
  assign T106 = T1310 ? 1'h0 : T107;
  assign T107 = T1308 ? reqDoneWire_19 : T108;
  assign T108 = T1288 ? 1'h0 : T109;
  assign T109 = T1286 ? reqDoneWire_19 : T110;
  assign T110 = T1266 ? 1'h0 : T111;
  assign T111 = T1264 ? reqDoneWire_19 : T112;
  assign T112 = T1244 ? 1'h0 : T113;
  assign T113 = T1242 ? reqDoneWire_19 : T114;
  assign T114 = T1222 ? 1'h0 : T115;
  assign T115 = T1220 ? reqDoneWire_19 : T116;
  assign T116 = T1200 ? 1'h0 : T117;
  assign T117 = T1198 ? reqDoneWire_19 : T118;
  assign T118 = T1178 ? 1'h0 : T119;
  assign T119 = T1176 ? reqDoneWire_19 : T120;
  assign T120 = T1156 ? 1'h0 : T121;
  assign T121 = T1154 ? reqDoneWire_19 : T122;
  assign T122 = T1134 ? 1'h0 : T123;
  assign T123 = T1132 ? reqDoneWire_19 : T124;
  assign T124 = T1112 ? 1'h0 : T125;
  assign T125 = T1110 ? reqDoneWire_19 : T126;
  assign T126 = T1090 ? 1'h0 : T127;
  assign T127 = T1088 ? reqDoneWire_19 : T128;
  assign T128 = T1068 ? 1'h0 : T129;
  assign T129 = T1066 ? reqDoneWire_19 : T130;
  assign T130 = T86 ? 1'h0 : reqDone_19;
  assign T136 = computeEnable & T137;
  assign T137 = T132 ^ 1'h1;
  assign T138 = T189 & reqDoneWire_18;
  assign reqDoneWire_18 = T139;
  assign T139 = T187 ? reqDone_18 : T140;
  assign T140 = T182 ? 1'h1 : T141;
  assign T141 = computeEnable ? reqDone_18 : 1'h0;
  assign T182 = computeEnable & T183;
  assign T183 = nextRequest_18 | T184;
  assign T184 = ~ io_outLocValid_18;
  assign nextRequest_18 = T185;
  assign T185 = T186 ? 1'h0 : io_seqProceed_18;
  assign T186 = io_seqProceed_18 ^ 1'h1;
  assign T1658 = reset ? 1'h0 : T142;
  assign T142 = T1484 ? reqDoneWire_18 : T143;
  assign T143 = T1464 ? 1'h0 : T144;
  assign T144 = T1462 ? reqDoneWire_18 : T145;
  assign T145 = T1442 ? 1'h0 : T146;
  assign T146 = T1440 ? reqDoneWire_18 : T147;
  assign T147 = T1420 ? 1'h0 : T148;
  assign T148 = T1418 ? reqDoneWire_18 : T149;
  assign T149 = T1398 ? 1'h0 : T150;
  assign T150 = T1396 ? reqDoneWire_18 : T151;
  assign T151 = T1376 ? 1'h0 : T152;
  assign T152 = T1374 ? reqDoneWire_18 : T153;
  assign T153 = T1354 ? 1'h0 : T154;
  assign T154 = T1352 ? reqDoneWire_18 : T155;
  assign T155 = T1332 ? 1'h0 : T156;
  assign T156 = T1330 ? reqDoneWire_18 : T157;
  assign T157 = T1310 ? 1'h0 : T158;
  assign T158 = T1308 ? reqDoneWire_18 : T159;
  assign T159 = T1288 ? 1'h0 : T160;
  assign T160 = T1286 ? reqDoneWire_18 : T161;
  assign T161 = T1266 ? 1'h0 : T162;
  assign T162 = T1264 ? reqDoneWire_18 : T163;
  assign T163 = T1244 ? 1'h0 : T164;
  assign T164 = T1242 ? reqDoneWire_18 : T165;
  assign T165 = T1222 ? 1'h0 : T166;
  assign T166 = T1220 ? reqDoneWire_18 : T167;
  assign T167 = T1200 ? 1'h0 : T168;
  assign T168 = T1198 ? reqDoneWire_18 : T169;
  assign T169 = T1178 ? 1'h0 : T170;
  assign T170 = T1176 ? reqDoneWire_18 : T171;
  assign T171 = T1156 ? 1'h0 : T172;
  assign T172 = T1154 ? reqDoneWire_18 : T173;
  assign T173 = T1134 ? 1'h0 : T174;
  assign T174 = T1132 ? reqDoneWire_18 : T175;
  assign T175 = T1112 ? 1'h0 : T176;
  assign T176 = T1110 ? reqDoneWire_18 : T177;
  assign T177 = T1090 ? 1'h0 : T178;
  assign T178 = T1088 ? reqDoneWire_18 : T179;
  assign T179 = T1068 ? 1'h0 : T180;
  assign T180 = T1066 ? reqDoneWire_18 : T181;
  assign T181 = T86 ? 1'h0 : reqDone_18;
  assign T187 = computeEnable & T188;
  assign T188 = T183 ^ 1'h1;
  assign T189 = T240 & reqDoneWire_17;
  assign reqDoneWire_17 = T190;
  assign T190 = T238 ? reqDone_17 : T191;
  assign T191 = T233 ? 1'h1 : T192;
  assign T192 = computeEnable ? reqDone_17 : 1'h0;
  assign T233 = computeEnable & T234;
  assign T234 = nextRequest_17 | T235;
  assign T235 = ~ io_outLocValid_17;
  assign nextRequest_17 = T236;
  assign T236 = T237 ? 1'h0 : io_seqProceed_17;
  assign T237 = io_seqProceed_17 ^ 1'h1;
  assign T1659 = reset ? 1'h0 : T193;
  assign T193 = T1484 ? reqDoneWire_17 : T194;
  assign T194 = T1464 ? 1'h0 : T195;
  assign T195 = T1462 ? reqDoneWire_17 : T196;
  assign T196 = T1442 ? 1'h0 : T197;
  assign T197 = T1440 ? reqDoneWire_17 : T198;
  assign T198 = T1420 ? 1'h0 : T199;
  assign T199 = T1418 ? reqDoneWire_17 : T200;
  assign T200 = T1398 ? 1'h0 : T201;
  assign T201 = T1396 ? reqDoneWire_17 : T202;
  assign T202 = T1376 ? 1'h0 : T203;
  assign T203 = T1374 ? reqDoneWire_17 : T204;
  assign T204 = T1354 ? 1'h0 : T205;
  assign T205 = T1352 ? reqDoneWire_17 : T206;
  assign T206 = T1332 ? 1'h0 : T207;
  assign T207 = T1330 ? reqDoneWire_17 : T208;
  assign T208 = T1310 ? 1'h0 : T209;
  assign T209 = T1308 ? reqDoneWire_17 : T210;
  assign T210 = T1288 ? 1'h0 : T211;
  assign T211 = T1286 ? reqDoneWire_17 : T212;
  assign T212 = T1266 ? 1'h0 : T213;
  assign T213 = T1264 ? reqDoneWire_17 : T214;
  assign T214 = T1244 ? 1'h0 : T215;
  assign T215 = T1242 ? reqDoneWire_17 : T216;
  assign T216 = T1222 ? 1'h0 : T217;
  assign T217 = T1220 ? reqDoneWire_17 : T218;
  assign T218 = T1200 ? 1'h0 : T219;
  assign T219 = T1198 ? reqDoneWire_17 : T220;
  assign T220 = T1178 ? 1'h0 : T221;
  assign T221 = T1176 ? reqDoneWire_17 : T222;
  assign T222 = T1156 ? 1'h0 : T223;
  assign T223 = T1154 ? reqDoneWire_17 : T224;
  assign T224 = T1134 ? 1'h0 : T225;
  assign T225 = T1132 ? reqDoneWire_17 : T226;
  assign T226 = T1112 ? 1'h0 : T227;
  assign T227 = T1110 ? reqDoneWire_17 : T228;
  assign T228 = T1090 ? 1'h0 : T229;
  assign T229 = T1088 ? reqDoneWire_17 : T230;
  assign T230 = T1068 ? 1'h0 : T231;
  assign T231 = T1066 ? reqDoneWire_17 : T232;
  assign T232 = T86 ? 1'h0 : reqDone_17;
  assign T238 = computeEnable & T239;
  assign T239 = T234 ^ 1'h1;
  assign T240 = T291 & reqDoneWire_16;
  assign reqDoneWire_16 = T241;
  assign T241 = T289 ? reqDone_16 : T242;
  assign T242 = T284 ? 1'h1 : T243;
  assign T243 = computeEnable ? reqDone_16 : 1'h0;
  assign T284 = computeEnable & T285;
  assign T285 = nextRequest_16 | T286;
  assign T286 = ~ io_outLocValid_16;
  assign nextRequest_16 = T287;
  assign T287 = T288 ? 1'h0 : io_seqProceed_16;
  assign T288 = io_seqProceed_16 ^ 1'h1;
  assign T1660 = reset ? 1'h0 : T244;
  assign T244 = T1484 ? reqDoneWire_16 : T245;
  assign T245 = T1464 ? 1'h0 : T246;
  assign T246 = T1462 ? reqDoneWire_16 : T247;
  assign T247 = T1442 ? 1'h0 : T248;
  assign T248 = T1440 ? reqDoneWire_16 : T249;
  assign T249 = T1420 ? 1'h0 : T250;
  assign T250 = T1418 ? reqDoneWire_16 : T251;
  assign T251 = T1398 ? 1'h0 : T252;
  assign T252 = T1396 ? reqDoneWire_16 : T253;
  assign T253 = T1376 ? 1'h0 : T254;
  assign T254 = T1374 ? reqDoneWire_16 : T255;
  assign T255 = T1354 ? 1'h0 : T256;
  assign T256 = T1352 ? reqDoneWire_16 : T257;
  assign T257 = T1332 ? 1'h0 : T258;
  assign T258 = T1330 ? reqDoneWire_16 : T259;
  assign T259 = T1310 ? 1'h0 : T260;
  assign T260 = T1308 ? reqDoneWire_16 : T261;
  assign T261 = T1288 ? 1'h0 : T262;
  assign T262 = T1286 ? reqDoneWire_16 : T263;
  assign T263 = T1266 ? 1'h0 : T264;
  assign T264 = T1264 ? reqDoneWire_16 : T265;
  assign T265 = T1244 ? 1'h0 : T266;
  assign T266 = T1242 ? reqDoneWire_16 : T267;
  assign T267 = T1222 ? 1'h0 : T268;
  assign T268 = T1220 ? reqDoneWire_16 : T269;
  assign T269 = T1200 ? 1'h0 : T270;
  assign T270 = T1198 ? reqDoneWire_16 : T271;
  assign T271 = T1178 ? 1'h0 : T272;
  assign T272 = T1176 ? reqDoneWire_16 : T273;
  assign T273 = T1156 ? 1'h0 : T274;
  assign T274 = T1154 ? reqDoneWire_16 : T275;
  assign T275 = T1134 ? 1'h0 : T276;
  assign T276 = T1132 ? reqDoneWire_16 : T277;
  assign T277 = T1112 ? 1'h0 : T278;
  assign T278 = T1110 ? reqDoneWire_16 : T279;
  assign T279 = T1090 ? 1'h0 : T280;
  assign T280 = T1088 ? reqDoneWire_16 : T281;
  assign T281 = T1068 ? 1'h0 : T282;
  assign T282 = T1066 ? reqDoneWire_16 : T283;
  assign T283 = T86 ? 1'h0 : reqDone_16;
  assign T289 = computeEnable & T290;
  assign T290 = T285 ^ 1'h1;
  assign T291 = T342 & reqDoneWire_15;
  assign reqDoneWire_15 = T292;
  assign T292 = T340 ? reqDone_15 : T293;
  assign T293 = T335 ? 1'h1 : T294;
  assign T294 = computeEnable ? reqDone_15 : 1'h0;
  assign T335 = computeEnable & T336;
  assign T336 = nextRequest_15 | T337;
  assign T337 = ~ io_outLocValid_15;
  assign nextRequest_15 = T338;
  assign T338 = T339 ? 1'h0 : io_seqProceed_15;
  assign T339 = io_seqProceed_15 ^ 1'h1;
  assign T1661 = reset ? 1'h0 : T295;
  assign T295 = T1484 ? reqDoneWire_15 : T296;
  assign T296 = T1464 ? 1'h0 : T297;
  assign T297 = T1462 ? reqDoneWire_15 : T298;
  assign T298 = T1442 ? 1'h0 : T299;
  assign T299 = T1440 ? reqDoneWire_15 : T300;
  assign T300 = T1420 ? 1'h0 : T301;
  assign T301 = T1418 ? reqDoneWire_15 : T302;
  assign T302 = T1398 ? 1'h0 : T303;
  assign T303 = T1396 ? reqDoneWire_15 : T304;
  assign T304 = T1376 ? 1'h0 : T305;
  assign T305 = T1374 ? reqDoneWire_15 : T306;
  assign T306 = T1354 ? 1'h0 : T307;
  assign T307 = T1352 ? reqDoneWire_15 : T308;
  assign T308 = T1332 ? 1'h0 : T309;
  assign T309 = T1330 ? reqDoneWire_15 : T310;
  assign T310 = T1310 ? 1'h0 : T311;
  assign T311 = T1308 ? reqDoneWire_15 : T312;
  assign T312 = T1288 ? 1'h0 : T313;
  assign T313 = T1286 ? reqDoneWire_15 : T314;
  assign T314 = T1266 ? 1'h0 : T315;
  assign T315 = T1264 ? reqDoneWire_15 : T316;
  assign T316 = T1244 ? 1'h0 : T317;
  assign T317 = T1242 ? reqDoneWire_15 : T318;
  assign T318 = T1222 ? 1'h0 : T319;
  assign T319 = T1220 ? reqDoneWire_15 : T320;
  assign T320 = T1200 ? 1'h0 : T321;
  assign T321 = T1198 ? reqDoneWire_15 : T322;
  assign T322 = T1178 ? 1'h0 : T323;
  assign T323 = T1176 ? reqDoneWire_15 : T324;
  assign T324 = T1156 ? 1'h0 : T325;
  assign T325 = T1154 ? reqDoneWire_15 : T326;
  assign T326 = T1134 ? 1'h0 : T327;
  assign T327 = T1132 ? reqDoneWire_15 : T328;
  assign T328 = T1112 ? 1'h0 : T329;
  assign T329 = T1110 ? reqDoneWire_15 : T330;
  assign T330 = T1090 ? 1'h0 : T331;
  assign T331 = T1088 ? reqDoneWire_15 : T332;
  assign T332 = T1068 ? 1'h0 : T333;
  assign T333 = T1066 ? reqDoneWire_15 : T334;
  assign T334 = T86 ? 1'h0 : reqDone_15;
  assign T340 = computeEnable & T341;
  assign T341 = T336 ^ 1'h1;
  assign T342 = T393 & reqDoneWire_14;
  assign reqDoneWire_14 = T343;
  assign T343 = T391 ? reqDone_14 : T344;
  assign T344 = T386 ? 1'h1 : T345;
  assign T345 = computeEnable ? reqDone_14 : 1'h0;
  assign T386 = computeEnable & T387;
  assign T387 = nextRequest_14 | T388;
  assign T388 = ~ io_outLocValid_14;
  assign nextRequest_14 = T389;
  assign T389 = T390 ? 1'h0 : io_seqProceed_14;
  assign T390 = io_seqProceed_14 ^ 1'h1;
  assign T1662 = reset ? 1'h0 : T346;
  assign T346 = T1484 ? reqDoneWire_14 : T347;
  assign T347 = T1464 ? 1'h0 : T348;
  assign T348 = T1462 ? reqDoneWire_14 : T349;
  assign T349 = T1442 ? 1'h0 : T350;
  assign T350 = T1440 ? reqDoneWire_14 : T351;
  assign T351 = T1420 ? 1'h0 : T352;
  assign T352 = T1418 ? reqDoneWire_14 : T353;
  assign T353 = T1398 ? 1'h0 : T354;
  assign T354 = T1396 ? reqDoneWire_14 : T355;
  assign T355 = T1376 ? 1'h0 : T356;
  assign T356 = T1374 ? reqDoneWire_14 : T357;
  assign T357 = T1354 ? 1'h0 : T358;
  assign T358 = T1352 ? reqDoneWire_14 : T359;
  assign T359 = T1332 ? 1'h0 : T360;
  assign T360 = T1330 ? reqDoneWire_14 : T361;
  assign T361 = T1310 ? 1'h0 : T362;
  assign T362 = T1308 ? reqDoneWire_14 : T363;
  assign T363 = T1288 ? 1'h0 : T364;
  assign T364 = T1286 ? reqDoneWire_14 : T365;
  assign T365 = T1266 ? 1'h0 : T366;
  assign T366 = T1264 ? reqDoneWire_14 : T367;
  assign T367 = T1244 ? 1'h0 : T368;
  assign T368 = T1242 ? reqDoneWire_14 : T369;
  assign T369 = T1222 ? 1'h0 : T370;
  assign T370 = T1220 ? reqDoneWire_14 : T371;
  assign T371 = T1200 ? 1'h0 : T372;
  assign T372 = T1198 ? reqDoneWire_14 : T373;
  assign T373 = T1178 ? 1'h0 : T374;
  assign T374 = T1176 ? reqDoneWire_14 : T375;
  assign T375 = T1156 ? 1'h0 : T376;
  assign T376 = T1154 ? reqDoneWire_14 : T377;
  assign T377 = T1134 ? 1'h0 : T378;
  assign T378 = T1132 ? reqDoneWire_14 : T379;
  assign T379 = T1112 ? 1'h0 : T380;
  assign T380 = T1110 ? reqDoneWire_14 : T381;
  assign T381 = T1090 ? 1'h0 : T382;
  assign T382 = T1088 ? reqDoneWire_14 : T383;
  assign T383 = T1068 ? 1'h0 : T384;
  assign T384 = T1066 ? reqDoneWire_14 : T385;
  assign T385 = T86 ? 1'h0 : reqDone_14;
  assign T391 = computeEnable & T392;
  assign T392 = T387 ^ 1'h1;
  assign T393 = T444 & reqDoneWire_13;
  assign reqDoneWire_13 = T394;
  assign T394 = T442 ? reqDone_13 : T395;
  assign T395 = T437 ? 1'h1 : T396;
  assign T396 = computeEnable ? reqDone_13 : 1'h0;
  assign T437 = computeEnable & T438;
  assign T438 = nextRequest_13 | T439;
  assign T439 = ~ io_outLocValid_13;
  assign nextRequest_13 = T440;
  assign T440 = T441 ? 1'h0 : io_seqProceed_13;
  assign T441 = io_seqProceed_13 ^ 1'h1;
  assign T1663 = reset ? 1'h0 : T397;
  assign T397 = T1484 ? reqDoneWire_13 : T398;
  assign T398 = T1464 ? 1'h0 : T399;
  assign T399 = T1462 ? reqDoneWire_13 : T400;
  assign T400 = T1442 ? 1'h0 : T401;
  assign T401 = T1440 ? reqDoneWire_13 : T402;
  assign T402 = T1420 ? 1'h0 : T403;
  assign T403 = T1418 ? reqDoneWire_13 : T404;
  assign T404 = T1398 ? 1'h0 : T405;
  assign T405 = T1396 ? reqDoneWire_13 : T406;
  assign T406 = T1376 ? 1'h0 : T407;
  assign T407 = T1374 ? reqDoneWire_13 : T408;
  assign T408 = T1354 ? 1'h0 : T409;
  assign T409 = T1352 ? reqDoneWire_13 : T410;
  assign T410 = T1332 ? 1'h0 : T411;
  assign T411 = T1330 ? reqDoneWire_13 : T412;
  assign T412 = T1310 ? 1'h0 : T413;
  assign T413 = T1308 ? reqDoneWire_13 : T414;
  assign T414 = T1288 ? 1'h0 : T415;
  assign T415 = T1286 ? reqDoneWire_13 : T416;
  assign T416 = T1266 ? 1'h0 : T417;
  assign T417 = T1264 ? reqDoneWire_13 : T418;
  assign T418 = T1244 ? 1'h0 : T419;
  assign T419 = T1242 ? reqDoneWire_13 : T420;
  assign T420 = T1222 ? 1'h0 : T421;
  assign T421 = T1220 ? reqDoneWire_13 : T422;
  assign T422 = T1200 ? 1'h0 : T423;
  assign T423 = T1198 ? reqDoneWire_13 : T424;
  assign T424 = T1178 ? 1'h0 : T425;
  assign T425 = T1176 ? reqDoneWire_13 : T426;
  assign T426 = T1156 ? 1'h0 : T427;
  assign T427 = T1154 ? reqDoneWire_13 : T428;
  assign T428 = T1134 ? 1'h0 : T429;
  assign T429 = T1132 ? reqDoneWire_13 : T430;
  assign T430 = T1112 ? 1'h0 : T431;
  assign T431 = T1110 ? reqDoneWire_13 : T432;
  assign T432 = T1090 ? 1'h0 : T433;
  assign T433 = T1088 ? reqDoneWire_13 : T434;
  assign T434 = T1068 ? 1'h0 : T435;
  assign T435 = T1066 ? reqDoneWire_13 : T436;
  assign T436 = T86 ? 1'h0 : reqDone_13;
  assign T442 = computeEnable & T443;
  assign T443 = T438 ^ 1'h1;
  assign T444 = T495 & reqDoneWire_12;
  assign reqDoneWire_12 = T445;
  assign T445 = T493 ? reqDone_12 : T446;
  assign T446 = T488 ? 1'h1 : T447;
  assign T447 = computeEnable ? reqDone_12 : 1'h0;
  assign T488 = computeEnable & T489;
  assign T489 = nextRequest_12 | T490;
  assign T490 = ~ io_outLocValid_12;
  assign nextRequest_12 = T491;
  assign T491 = T492 ? 1'h0 : io_seqProceed_12;
  assign T492 = io_seqProceed_12 ^ 1'h1;
  assign T1664 = reset ? 1'h0 : T448;
  assign T448 = T1484 ? reqDoneWire_12 : T449;
  assign T449 = T1464 ? 1'h0 : T450;
  assign T450 = T1462 ? reqDoneWire_12 : T451;
  assign T451 = T1442 ? 1'h0 : T452;
  assign T452 = T1440 ? reqDoneWire_12 : T453;
  assign T453 = T1420 ? 1'h0 : T454;
  assign T454 = T1418 ? reqDoneWire_12 : T455;
  assign T455 = T1398 ? 1'h0 : T456;
  assign T456 = T1396 ? reqDoneWire_12 : T457;
  assign T457 = T1376 ? 1'h0 : T458;
  assign T458 = T1374 ? reqDoneWire_12 : T459;
  assign T459 = T1354 ? 1'h0 : T460;
  assign T460 = T1352 ? reqDoneWire_12 : T461;
  assign T461 = T1332 ? 1'h0 : T462;
  assign T462 = T1330 ? reqDoneWire_12 : T463;
  assign T463 = T1310 ? 1'h0 : T464;
  assign T464 = T1308 ? reqDoneWire_12 : T465;
  assign T465 = T1288 ? 1'h0 : T466;
  assign T466 = T1286 ? reqDoneWire_12 : T467;
  assign T467 = T1266 ? 1'h0 : T468;
  assign T468 = T1264 ? reqDoneWire_12 : T469;
  assign T469 = T1244 ? 1'h0 : T470;
  assign T470 = T1242 ? reqDoneWire_12 : T471;
  assign T471 = T1222 ? 1'h0 : T472;
  assign T472 = T1220 ? reqDoneWire_12 : T473;
  assign T473 = T1200 ? 1'h0 : T474;
  assign T474 = T1198 ? reqDoneWire_12 : T475;
  assign T475 = T1178 ? 1'h0 : T476;
  assign T476 = T1176 ? reqDoneWire_12 : T477;
  assign T477 = T1156 ? 1'h0 : T478;
  assign T478 = T1154 ? reqDoneWire_12 : T479;
  assign T479 = T1134 ? 1'h0 : T480;
  assign T480 = T1132 ? reqDoneWire_12 : T481;
  assign T481 = T1112 ? 1'h0 : T482;
  assign T482 = T1110 ? reqDoneWire_12 : T483;
  assign T483 = T1090 ? 1'h0 : T484;
  assign T484 = T1088 ? reqDoneWire_12 : T485;
  assign T485 = T1068 ? 1'h0 : T486;
  assign T486 = T1066 ? reqDoneWire_12 : T487;
  assign T487 = T86 ? 1'h0 : reqDone_12;
  assign T493 = computeEnable & T494;
  assign T494 = T489 ^ 1'h1;
  assign T495 = T546 & reqDoneWire_11;
  assign reqDoneWire_11 = T496;
  assign T496 = T544 ? reqDone_11 : T497;
  assign T497 = T539 ? 1'h1 : T498;
  assign T498 = computeEnable ? reqDone_11 : 1'h0;
  assign T539 = computeEnable & T540;
  assign T540 = nextRequest_11 | T541;
  assign T541 = ~ io_outLocValid_11;
  assign nextRequest_11 = T542;
  assign T542 = T543 ? 1'h0 : io_seqProceed_11;
  assign T543 = io_seqProceed_11 ^ 1'h1;
  assign T1665 = reset ? 1'h0 : T499;
  assign T499 = T1484 ? reqDoneWire_11 : T500;
  assign T500 = T1464 ? 1'h0 : T501;
  assign T501 = T1462 ? reqDoneWire_11 : T502;
  assign T502 = T1442 ? 1'h0 : T503;
  assign T503 = T1440 ? reqDoneWire_11 : T504;
  assign T504 = T1420 ? 1'h0 : T505;
  assign T505 = T1418 ? reqDoneWire_11 : T506;
  assign T506 = T1398 ? 1'h0 : T507;
  assign T507 = T1396 ? reqDoneWire_11 : T508;
  assign T508 = T1376 ? 1'h0 : T509;
  assign T509 = T1374 ? reqDoneWire_11 : T510;
  assign T510 = T1354 ? 1'h0 : T511;
  assign T511 = T1352 ? reqDoneWire_11 : T512;
  assign T512 = T1332 ? 1'h0 : T513;
  assign T513 = T1330 ? reqDoneWire_11 : T514;
  assign T514 = T1310 ? 1'h0 : T515;
  assign T515 = T1308 ? reqDoneWire_11 : T516;
  assign T516 = T1288 ? 1'h0 : T517;
  assign T517 = T1286 ? reqDoneWire_11 : T518;
  assign T518 = T1266 ? 1'h0 : T519;
  assign T519 = T1264 ? reqDoneWire_11 : T520;
  assign T520 = T1244 ? 1'h0 : T521;
  assign T521 = T1242 ? reqDoneWire_11 : T522;
  assign T522 = T1222 ? 1'h0 : T523;
  assign T523 = T1220 ? reqDoneWire_11 : T524;
  assign T524 = T1200 ? 1'h0 : T525;
  assign T525 = T1198 ? reqDoneWire_11 : T526;
  assign T526 = T1178 ? 1'h0 : T527;
  assign T527 = T1176 ? reqDoneWire_11 : T528;
  assign T528 = T1156 ? 1'h0 : T529;
  assign T529 = T1154 ? reqDoneWire_11 : T530;
  assign T530 = T1134 ? 1'h0 : T531;
  assign T531 = T1132 ? reqDoneWire_11 : T532;
  assign T532 = T1112 ? 1'h0 : T533;
  assign T533 = T1110 ? reqDoneWire_11 : T534;
  assign T534 = T1090 ? 1'h0 : T535;
  assign T535 = T1088 ? reqDoneWire_11 : T536;
  assign T536 = T1068 ? 1'h0 : T537;
  assign T537 = T1066 ? reqDoneWire_11 : T538;
  assign T538 = T86 ? 1'h0 : reqDone_11;
  assign T544 = computeEnable & T545;
  assign T545 = T540 ^ 1'h1;
  assign T546 = T597 & reqDoneWire_10;
  assign reqDoneWire_10 = T547;
  assign T547 = T595 ? reqDone_10 : T548;
  assign T548 = T590 ? 1'h1 : T549;
  assign T549 = computeEnable ? reqDone_10 : 1'h0;
  assign T590 = computeEnable & T591;
  assign T591 = nextRequest_10 | T592;
  assign T592 = ~ io_outLocValid_10;
  assign nextRequest_10 = T593;
  assign T593 = T594 ? 1'h0 : io_seqProceed_10;
  assign T594 = io_seqProceed_10 ^ 1'h1;
  assign T1666 = reset ? 1'h0 : T550;
  assign T550 = T1484 ? reqDoneWire_10 : T551;
  assign T551 = T1464 ? 1'h0 : T552;
  assign T552 = T1462 ? reqDoneWire_10 : T553;
  assign T553 = T1442 ? 1'h0 : T554;
  assign T554 = T1440 ? reqDoneWire_10 : T555;
  assign T555 = T1420 ? 1'h0 : T556;
  assign T556 = T1418 ? reqDoneWire_10 : T557;
  assign T557 = T1398 ? 1'h0 : T558;
  assign T558 = T1396 ? reqDoneWire_10 : T559;
  assign T559 = T1376 ? 1'h0 : T560;
  assign T560 = T1374 ? reqDoneWire_10 : T561;
  assign T561 = T1354 ? 1'h0 : T562;
  assign T562 = T1352 ? reqDoneWire_10 : T563;
  assign T563 = T1332 ? 1'h0 : T564;
  assign T564 = T1330 ? reqDoneWire_10 : T565;
  assign T565 = T1310 ? 1'h0 : T566;
  assign T566 = T1308 ? reqDoneWire_10 : T567;
  assign T567 = T1288 ? 1'h0 : T568;
  assign T568 = T1286 ? reqDoneWire_10 : T569;
  assign T569 = T1266 ? 1'h0 : T570;
  assign T570 = T1264 ? reqDoneWire_10 : T571;
  assign T571 = T1244 ? 1'h0 : T572;
  assign T572 = T1242 ? reqDoneWire_10 : T573;
  assign T573 = T1222 ? 1'h0 : T574;
  assign T574 = T1220 ? reqDoneWire_10 : T575;
  assign T575 = T1200 ? 1'h0 : T576;
  assign T576 = T1198 ? reqDoneWire_10 : T577;
  assign T577 = T1178 ? 1'h0 : T578;
  assign T578 = T1176 ? reqDoneWire_10 : T579;
  assign T579 = T1156 ? 1'h0 : T580;
  assign T580 = T1154 ? reqDoneWire_10 : T581;
  assign T581 = T1134 ? 1'h0 : T582;
  assign T582 = T1132 ? reqDoneWire_10 : T583;
  assign T583 = T1112 ? 1'h0 : T584;
  assign T584 = T1110 ? reqDoneWire_10 : T585;
  assign T585 = T1090 ? 1'h0 : T586;
  assign T586 = T1088 ? reqDoneWire_10 : T587;
  assign T587 = T1068 ? 1'h0 : T588;
  assign T588 = T1066 ? reqDoneWire_10 : T589;
  assign T589 = T86 ? 1'h0 : reqDone_10;
  assign T595 = computeEnable & T596;
  assign T596 = T591 ^ 1'h1;
  assign T597 = T648 & reqDoneWire_9;
  assign reqDoneWire_9 = T598;
  assign T598 = T646 ? reqDone_9 : T599;
  assign T599 = T641 ? 1'h1 : T600;
  assign T600 = computeEnable ? reqDone_9 : 1'h0;
  assign T641 = computeEnable & T642;
  assign T642 = nextRequest_9 | T643;
  assign T643 = ~ io_outLocValid_9;
  assign nextRequest_9 = T644;
  assign T644 = T645 ? 1'h0 : io_seqProceed_9;
  assign T645 = io_seqProceed_9 ^ 1'h1;
  assign T1667 = reset ? 1'h0 : T601;
  assign T601 = T1484 ? reqDoneWire_9 : T602;
  assign T602 = T1464 ? 1'h0 : T603;
  assign T603 = T1462 ? reqDoneWire_9 : T604;
  assign T604 = T1442 ? 1'h0 : T605;
  assign T605 = T1440 ? reqDoneWire_9 : T606;
  assign T606 = T1420 ? 1'h0 : T607;
  assign T607 = T1418 ? reqDoneWire_9 : T608;
  assign T608 = T1398 ? 1'h0 : T609;
  assign T609 = T1396 ? reqDoneWire_9 : T610;
  assign T610 = T1376 ? 1'h0 : T611;
  assign T611 = T1374 ? reqDoneWire_9 : T612;
  assign T612 = T1354 ? 1'h0 : T613;
  assign T613 = T1352 ? reqDoneWire_9 : T614;
  assign T614 = T1332 ? 1'h0 : T615;
  assign T615 = T1330 ? reqDoneWire_9 : T616;
  assign T616 = T1310 ? 1'h0 : T617;
  assign T617 = T1308 ? reqDoneWire_9 : T618;
  assign T618 = T1288 ? 1'h0 : T619;
  assign T619 = T1286 ? reqDoneWire_9 : T620;
  assign T620 = T1266 ? 1'h0 : T621;
  assign T621 = T1264 ? reqDoneWire_9 : T622;
  assign T622 = T1244 ? 1'h0 : T623;
  assign T623 = T1242 ? reqDoneWire_9 : T624;
  assign T624 = T1222 ? 1'h0 : T625;
  assign T625 = T1220 ? reqDoneWire_9 : T626;
  assign T626 = T1200 ? 1'h0 : T627;
  assign T627 = T1198 ? reqDoneWire_9 : T628;
  assign T628 = T1178 ? 1'h0 : T629;
  assign T629 = T1176 ? reqDoneWire_9 : T630;
  assign T630 = T1156 ? 1'h0 : T631;
  assign T631 = T1154 ? reqDoneWire_9 : T632;
  assign T632 = T1134 ? 1'h0 : T633;
  assign T633 = T1132 ? reqDoneWire_9 : T634;
  assign T634 = T1112 ? 1'h0 : T635;
  assign T635 = T1110 ? reqDoneWire_9 : T636;
  assign T636 = T1090 ? 1'h0 : T637;
  assign T637 = T1088 ? reqDoneWire_9 : T638;
  assign T638 = T1068 ? 1'h0 : T639;
  assign T639 = T1066 ? reqDoneWire_9 : T640;
  assign T640 = T86 ? 1'h0 : reqDone_9;
  assign T646 = computeEnable & T647;
  assign T647 = T642 ^ 1'h1;
  assign T648 = T699 & reqDoneWire_8;
  assign reqDoneWire_8 = T649;
  assign T649 = T697 ? reqDone_8 : T650;
  assign T650 = T692 ? 1'h1 : T651;
  assign T651 = computeEnable ? reqDone_8 : 1'h0;
  assign T692 = computeEnable & T693;
  assign T693 = nextRequest_8 | T694;
  assign T694 = ~ io_outLocValid_8;
  assign nextRequest_8 = T695;
  assign T695 = T696 ? 1'h0 : io_seqProceed_8;
  assign T696 = io_seqProceed_8 ^ 1'h1;
  assign T1668 = reset ? 1'h0 : T652;
  assign T652 = T1484 ? reqDoneWire_8 : T653;
  assign T653 = T1464 ? 1'h0 : T654;
  assign T654 = T1462 ? reqDoneWire_8 : T655;
  assign T655 = T1442 ? 1'h0 : T656;
  assign T656 = T1440 ? reqDoneWire_8 : T657;
  assign T657 = T1420 ? 1'h0 : T658;
  assign T658 = T1418 ? reqDoneWire_8 : T659;
  assign T659 = T1398 ? 1'h0 : T660;
  assign T660 = T1396 ? reqDoneWire_8 : T661;
  assign T661 = T1376 ? 1'h0 : T662;
  assign T662 = T1374 ? reqDoneWire_8 : T663;
  assign T663 = T1354 ? 1'h0 : T664;
  assign T664 = T1352 ? reqDoneWire_8 : T665;
  assign T665 = T1332 ? 1'h0 : T666;
  assign T666 = T1330 ? reqDoneWire_8 : T667;
  assign T667 = T1310 ? 1'h0 : T668;
  assign T668 = T1308 ? reqDoneWire_8 : T669;
  assign T669 = T1288 ? 1'h0 : T670;
  assign T670 = T1286 ? reqDoneWire_8 : T671;
  assign T671 = T1266 ? 1'h0 : T672;
  assign T672 = T1264 ? reqDoneWire_8 : T673;
  assign T673 = T1244 ? 1'h0 : T674;
  assign T674 = T1242 ? reqDoneWire_8 : T675;
  assign T675 = T1222 ? 1'h0 : T676;
  assign T676 = T1220 ? reqDoneWire_8 : T677;
  assign T677 = T1200 ? 1'h0 : T678;
  assign T678 = T1198 ? reqDoneWire_8 : T679;
  assign T679 = T1178 ? 1'h0 : T680;
  assign T680 = T1176 ? reqDoneWire_8 : T681;
  assign T681 = T1156 ? 1'h0 : T682;
  assign T682 = T1154 ? reqDoneWire_8 : T683;
  assign T683 = T1134 ? 1'h0 : T684;
  assign T684 = T1132 ? reqDoneWire_8 : T685;
  assign T685 = T1112 ? 1'h0 : T686;
  assign T686 = T1110 ? reqDoneWire_8 : T687;
  assign T687 = T1090 ? 1'h0 : T688;
  assign T688 = T1088 ? reqDoneWire_8 : T689;
  assign T689 = T1068 ? 1'h0 : T690;
  assign T690 = T1066 ? reqDoneWire_8 : T691;
  assign T691 = T86 ? 1'h0 : reqDone_8;
  assign T697 = computeEnable & T698;
  assign T698 = T693 ^ 1'h1;
  assign T699 = T750 & reqDoneWire_7;
  assign reqDoneWire_7 = T700;
  assign T700 = T748 ? reqDone_7 : T701;
  assign T701 = T743 ? 1'h1 : T702;
  assign T702 = computeEnable ? reqDone_7 : 1'h0;
  assign T743 = computeEnable & T744;
  assign T744 = nextRequest_7 | T745;
  assign T745 = ~ io_outLocValid_7;
  assign nextRequest_7 = T746;
  assign T746 = T747 ? 1'h0 : io_seqProceed_7;
  assign T747 = io_seqProceed_7 ^ 1'h1;
  assign T1669 = reset ? 1'h0 : T703;
  assign T703 = T1484 ? reqDoneWire_7 : T704;
  assign T704 = T1464 ? 1'h0 : T705;
  assign T705 = T1462 ? reqDoneWire_7 : T706;
  assign T706 = T1442 ? 1'h0 : T707;
  assign T707 = T1440 ? reqDoneWire_7 : T708;
  assign T708 = T1420 ? 1'h0 : T709;
  assign T709 = T1418 ? reqDoneWire_7 : T710;
  assign T710 = T1398 ? 1'h0 : T711;
  assign T711 = T1396 ? reqDoneWire_7 : T712;
  assign T712 = T1376 ? 1'h0 : T713;
  assign T713 = T1374 ? reqDoneWire_7 : T714;
  assign T714 = T1354 ? 1'h0 : T715;
  assign T715 = T1352 ? reqDoneWire_7 : T716;
  assign T716 = T1332 ? 1'h0 : T717;
  assign T717 = T1330 ? reqDoneWire_7 : T718;
  assign T718 = T1310 ? 1'h0 : T719;
  assign T719 = T1308 ? reqDoneWire_7 : T720;
  assign T720 = T1288 ? 1'h0 : T721;
  assign T721 = T1286 ? reqDoneWire_7 : T722;
  assign T722 = T1266 ? 1'h0 : T723;
  assign T723 = T1264 ? reqDoneWire_7 : T724;
  assign T724 = T1244 ? 1'h0 : T725;
  assign T725 = T1242 ? reqDoneWire_7 : T726;
  assign T726 = T1222 ? 1'h0 : T727;
  assign T727 = T1220 ? reqDoneWire_7 : T728;
  assign T728 = T1200 ? 1'h0 : T729;
  assign T729 = T1198 ? reqDoneWire_7 : T730;
  assign T730 = T1178 ? 1'h0 : T731;
  assign T731 = T1176 ? reqDoneWire_7 : T732;
  assign T732 = T1156 ? 1'h0 : T733;
  assign T733 = T1154 ? reqDoneWire_7 : T734;
  assign T734 = T1134 ? 1'h0 : T735;
  assign T735 = T1132 ? reqDoneWire_7 : T736;
  assign T736 = T1112 ? 1'h0 : T737;
  assign T737 = T1110 ? reqDoneWire_7 : T738;
  assign T738 = T1090 ? 1'h0 : T739;
  assign T739 = T1088 ? reqDoneWire_7 : T740;
  assign T740 = T1068 ? 1'h0 : T741;
  assign T741 = T1066 ? reqDoneWire_7 : T742;
  assign T742 = T86 ? 1'h0 : reqDone_7;
  assign T748 = computeEnable & T749;
  assign T749 = T744 ^ 1'h1;
  assign T750 = T801 & reqDoneWire_6;
  assign reqDoneWire_6 = T751;
  assign T751 = T799 ? reqDone_6 : T752;
  assign T752 = T794 ? 1'h1 : T753;
  assign T753 = computeEnable ? reqDone_6 : 1'h0;
  assign T794 = computeEnable & T795;
  assign T795 = nextRequest_6 | T796;
  assign T796 = ~ io_outLocValid_6;
  assign nextRequest_6 = T797;
  assign T797 = T798 ? 1'h0 : io_seqProceed_6;
  assign T798 = io_seqProceed_6 ^ 1'h1;
  assign T1670 = reset ? 1'h0 : T754;
  assign T754 = T1484 ? reqDoneWire_6 : T755;
  assign T755 = T1464 ? 1'h0 : T756;
  assign T756 = T1462 ? reqDoneWire_6 : T757;
  assign T757 = T1442 ? 1'h0 : T758;
  assign T758 = T1440 ? reqDoneWire_6 : T759;
  assign T759 = T1420 ? 1'h0 : T760;
  assign T760 = T1418 ? reqDoneWire_6 : T761;
  assign T761 = T1398 ? 1'h0 : T762;
  assign T762 = T1396 ? reqDoneWire_6 : T763;
  assign T763 = T1376 ? 1'h0 : T764;
  assign T764 = T1374 ? reqDoneWire_6 : T765;
  assign T765 = T1354 ? 1'h0 : T766;
  assign T766 = T1352 ? reqDoneWire_6 : T767;
  assign T767 = T1332 ? 1'h0 : T768;
  assign T768 = T1330 ? reqDoneWire_6 : T769;
  assign T769 = T1310 ? 1'h0 : T770;
  assign T770 = T1308 ? reqDoneWire_6 : T771;
  assign T771 = T1288 ? 1'h0 : T772;
  assign T772 = T1286 ? reqDoneWire_6 : T773;
  assign T773 = T1266 ? 1'h0 : T774;
  assign T774 = T1264 ? reqDoneWire_6 : T775;
  assign T775 = T1244 ? 1'h0 : T776;
  assign T776 = T1242 ? reqDoneWire_6 : T777;
  assign T777 = T1222 ? 1'h0 : T778;
  assign T778 = T1220 ? reqDoneWire_6 : T779;
  assign T779 = T1200 ? 1'h0 : T780;
  assign T780 = T1198 ? reqDoneWire_6 : T781;
  assign T781 = T1178 ? 1'h0 : T782;
  assign T782 = T1176 ? reqDoneWire_6 : T783;
  assign T783 = T1156 ? 1'h0 : T784;
  assign T784 = T1154 ? reqDoneWire_6 : T785;
  assign T785 = T1134 ? 1'h0 : T786;
  assign T786 = T1132 ? reqDoneWire_6 : T787;
  assign T787 = T1112 ? 1'h0 : T788;
  assign T788 = T1110 ? reqDoneWire_6 : T789;
  assign T789 = T1090 ? 1'h0 : T790;
  assign T790 = T1088 ? reqDoneWire_6 : T791;
  assign T791 = T1068 ? 1'h0 : T792;
  assign T792 = T1066 ? reqDoneWire_6 : T793;
  assign T793 = T86 ? 1'h0 : reqDone_6;
  assign T799 = computeEnable & T800;
  assign T800 = T795 ^ 1'h1;
  assign T801 = T852 & reqDoneWire_5;
  assign reqDoneWire_5 = T802;
  assign T802 = T850 ? reqDone_5 : T803;
  assign T803 = T845 ? 1'h1 : T804;
  assign T804 = computeEnable ? reqDone_5 : 1'h0;
  assign T845 = computeEnable & T846;
  assign T846 = nextRequest_5 | T847;
  assign T847 = ~ io_outLocValid_5;
  assign nextRequest_5 = T848;
  assign T848 = T849 ? 1'h0 : io_seqProceed_5;
  assign T849 = io_seqProceed_5 ^ 1'h1;
  assign T1671 = reset ? 1'h0 : T805;
  assign T805 = T1484 ? reqDoneWire_5 : T806;
  assign T806 = T1464 ? 1'h0 : T807;
  assign T807 = T1462 ? reqDoneWire_5 : T808;
  assign T808 = T1442 ? 1'h0 : T809;
  assign T809 = T1440 ? reqDoneWire_5 : T810;
  assign T810 = T1420 ? 1'h0 : T811;
  assign T811 = T1418 ? reqDoneWire_5 : T812;
  assign T812 = T1398 ? 1'h0 : T813;
  assign T813 = T1396 ? reqDoneWire_5 : T814;
  assign T814 = T1376 ? 1'h0 : T815;
  assign T815 = T1374 ? reqDoneWire_5 : T816;
  assign T816 = T1354 ? 1'h0 : T817;
  assign T817 = T1352 ? reqDoneWire_5 : T818;
  assign T818 = T1332 ? 1'h0 : T819;
  assign T819 = T1330 ? reqDoneWire_5 : T820;
  assign T820 = T1310 ? 1'h0 : T821;
  assign T821 = T1308 ? reqDoneWire_5 : T822;
  assign T822 = T1288 ? 1'h0 : T823;
  assign T823 = T1286 ? reqDoneWire_5 : T824;
  assign T824 = T1266 ? 1'h0 : T825;
  assign T825 = T1264 ? reqDoneWire_5 : T826;
  assign T826 = T1244 ? 1'h0 : T827;
  assign T827 = T1242 ? reqDoneWire_5 : T828;
  assign T828 = T1222 ? 1'h0 : T829;
  assign T829 = T1220 ? reqDoneWire_5 : T830;
  assign T830 = T1200 ? 1'h0 : T831;
  assign T831 = T1198 ? reqDoneWire_5 : T832;
  assign T832 = T1178 ? 1'h0 : T833;
  assign T833 = T1176 ? reqDoneWire_5 : T834;
  assign T834 = T1156 ? 1'h0 : T835;
  assign T835 = T1154 ? reqDoneWire_5 : T836;
  assign T836 = T1134 ? 1'h0 : T837;
  assign T837 = T1132 ? reqDoneWire_5 : T838;
  assign T838 = T1112 ? 1'h0 : T839;
  assign T839 = T1110 ? reqDoneWire_5 : T840;
  assign T840 = T1090 ? 1'h0 : T841;
  assign T841 = T1088 ? reqDoneWire_5 : T842;
  assign T842 = T1068 ? 1'h0 : T843;
  assign T843 = T1066 ? reqDoneWire_5 : T844;
  assign T844 = T86 ? 1'h0 : reqDone_5;
  assign T850 = computeEnable & T851;
  assign T851 = T846 ^ 1'h1;
  assign T852 = T903 & reqDoneWire_4;
  assign reqDoneWire_4 = T853;
  assign T853 = T901 ? reqDone_4 : T854;
  assign T854 = T896 ? 1'h1 : T855;
  assign T855 = computeEnable ? reqDone_4 : 1'h0;
  assign T896 = computeEnable & T897;
  assign T897 = nextRequest_4 | T898;
  assign T898 = ~ io_outLocValid_4;
  assign nextRequest_4 = T899;
  assign T899 = T900 ? 1'h0 : io_seqProceed_4;
  assign T900 = io_seqProceed_4 ^ 1'h1;
  assign T1672 = reset ? 1'h0 : T856;
  assign T856 = T1484 ? reqDoneWire_4 : T857;
  assign T857 = T1464 ? 1'h0 : T858;
  assign T858 = T1462 ? reqDoneWire_4 : T859;
  assign T859 = T1442 ? 1'h0 : T860;
  assign T860 = T1440 ? reqDoneWire_4 : T861;
  assign T861 = T1420 ? 1'h0 : T862;
  assign T862 = T1418 ? reqDoneWire_4 : T863;
  assign T863 = T1398 ? 1'h0 : T864;
  assign T864 = T1396 ? reqDoneWire_4 : T865;
  assign T865 = T1376 ? 1'h0 : T866;
  assign T866 = T1374 ? reqDoneWire_4 : T867;
  assign T867 = T1354 ? 1'h0 : T868;
  assign T868 = T1352 ? reqDoneWire_4 : T869;
  assign T869 = T1332 ? 1'h0 : T870;
  assign T870 = T1330 ? reqDoneWire_4 : T871;
  assign T871 = T1310 ? 1'h0 : T872;
  assign T872 = T1308 ? reqDoneWire_4 : T873;
  assign T873 = T1288 ? 1'h0 : T874;
  assign T874 = T1286 ? reqDoneWire_4 : T875;
  assign T875 = T1266 ? 1'h0 : T876;
  assign T876 = T1264 ? reqDoneWire_4 : T877;
  assign T877 = T1244 ? 1'h0 : T878;
  assign T878 = T1242 ? reqDoneWire_4 : T879;
  assign T879 = T1222 ? 1'h0 : T880;
  assign T880 = T1220 ? reqDoneWire_4 : T881;
  assign T881 = T1200 ? 1'h0 : T882;
  assign T882 = T1198 ? reqDoneWire_4 : T883;
  assign T883 = T1178 ? 1'h0 : T884;
  assign T884 = T1176 ? reqDoneWire_4 : T885;
  assign T885 = T1156 ? 1'h0 : T886;
  assign T886 = T1154 ? reqDoneWire_4 : T887;
  assign T887 = T1134 ? 1'h0 : T888;
  assign T888 = T1132 ? reqDoneWire_4 : T889;
  assign T889 = T1112 ? 1'h0 : T890;
  assign T890 = T1110 ? reqDoneWire_4 : T891;
  assign T891 = T1090 ? 1'h0 : T892;
  assign T892 = T1088 ? reqDoneWire_4 : T893;
  assign T893 = T1068 ? 1'h0 : T894;
  assign T894 = T1066 ? reqDoneWire_4 : T895;
  assign T895 = T86 ? 1'h0 : reqDone_4;
  assign T901 = computeEnable & T902;
  assign T902 = T897 ^ 1'h1;
  assign T903 = T954 & reqDoneWire_3;
  assign reqDoneWire_3 = T904;
  assign T904 = T952 ? reqDone_3 : T905;
  assign T905 = T947 ? 1'h1 : T906;
  assign T906 = computeEnable ? reqDone_3 : 1'h0;
  assign T947 = computeEnable & T948;
  assign T948 = nextRequest_3 | T949;
  assign T949 = ~ io_outLocValid_3;
  assign nextRequest_3 = T950;
  assign T950 = T951 ? 1'h0 : io_seqProceed_3;
  assign T951 = io_seqProceed_3 ^ 1'h1;
  assign T1673 = reset ? 1'h0 : T907;
  assign T907 = T1484 ? reqDoneWire_3 : T908;
  assign T908 = T1464 ? 1'h0 : T909;
  assign T909 = T1462 ? reqDoneWire_3 : T910;
  assign T910 = T1442 ? 1'h0 : T911;
  assign T911 = T1440 ? reqDoneWire_3 : T912;
  assign T912 = T1420 ? 1'h0 : T913;
  assign T913 = T1418 ? reqDoneWire_3 : T914;
  assign T914 = T1398 ? 1'h0 : T915;
  assign T915 = T1396 ? reqDoneWire_3 : T916;
  assign T916 = T1376 ? 1'h0 : T917;
  assign T917 = T1374 ? reqDoneWire_3 : T918;
  assign T918 = T1354 ? 1'h0 : T919;
  assign T919 = T1352 ? reqDoneWire_3 : T920;
  assign T920 = T1332 ? 1'h0 : T921;
  assign T921 = T1330 ? reqDoneWire_3 : T922;
  assign T922 = T1310 ? 1'h0 : T923;
  assign T923 = T1308 ? reqDoneWire_3 : T924;
  assign T924 = T1288 ? 1'h0 : T925;
  assign T925 = T1286 ? reqDoneWire_3 : T926;
  assign T926 = T1266 ? 1'h0 : T927;
  assign T927 = T1264 ? reqDoneWire_3 : T928;
  assign T928 = T1244 ? 1'h0 : T929;
  assign T929 = T1242 ? reqDoneWire_3 : T930;
  assign T930 = T1222 ? 1'h0 : T931;
  assign T931 = T1220 ? reqDoneWire_3 : T932;
  assign T932 = T1200 ? 1'h0 : T933;
  assign T933 = T1198 ? reqDoneWire_3 : T934;
  assign T934 = T1178 ? 1'h0 : T935;
  assign T935 = T1176 ? reqDoneWire_3 : T936;
  assign T936 = T1156 ? 1'h0 : T937;
  assign T937 = T1154 ? reqDoneWire_3 : T938;
  assign T938 = T1134 ? 1'h0 : T939;
  assign T939 = T1132 ? reqDoneWire_3 : T940;
  assign T940 = T1112 ? 1'h0 : T941;
  assign T941 = T1110 ? reqDoneWire_3 : T942;
  assign T942 = T1090 ? 1'h0 : T943;
  assign T943 = T1088 ? reqDoneWire_3 : T944;
  assign T944 = T1068 ? 1'h0 : T945;
  assign T945 = T1066 ? reqDoneWire_3 : T946;
  assign T946 = T86 ? 1'h0 : reqDone_3;
  assign T952 = computeEnable & T953;
  assign T953 = T948 ^ 1'h1;
  assign T954 = T1005 & reqDoneWire_2;
  assign reqDoneWire_2 = T955;
  assign T955 = T1003 ? reqDone_2 : T956;
  assign T956 = T998 ? 1'h1 : T957;
  assign T957 = computeEnable ? reqDone_2 : 1'h0;
  assign T998 = computeEnable & T999;
  assign T999 = nextRequest_2 | T1000;
  assign T1000 = ~ io_outLocValid_2;
  assign nextRequest_2 = T1001;
  assign T1001 = T1002 ? 1'h0 : io_seqProceed_2;
  assign T1002 = io_seqProceed_2 ^ 1'h1;
  assign T1674 = reset ? 1'h0 : T958;
  assign T958 = T1484 ? reqDoneWire_2 : T959;
  assign T959 = T1464 ? 1'h0 : T960;
  assign T960 = T1462 ? reqDoneWire_2 : T961;
  assign T961 = T1442 ? 1'h0 : T962;
  assign T962 = T1440 ? reqDoneWire_2 : T963;
  assign T963 = T1420 ? 1'h0 : T964;
  assign T964 = T1418 ? reqDoneWire_2 : T965;
  assign T965 = T1398 ? 1'h0 : T966;
  assign T966 = T1396 ? reqDoneWire_2 : T967;
  assign T967 = T1376 ? 1'h0 : T968;
  assign T968 = T1374 ? reqDoneWire_2 : T969;
  assign T969 = T1354 ? 1'h0 : T970;
  assign T970 = T1352 ? reqDoneWire_2 : T971;
  assign T971 = T1332 ? 1'h0 : T972;
  assign T972 = T1330 ? reqDoneWire_2 : T973;
  assign T973 = T1310 ? 1'h0 : T974;
  assign T974 = T1308 ? reqDoneWire_2 : T975;
  assign T975 = T1288 ? 1'h0 : T976;
  assign T976 = T1286 ? reqDoneWire_2 : T977;
  assign T977 = T1266 ? 1'h0 : T978;
  assign T978 = T1264 ? reqDoneWire_2 : T979;
  assign T979 = T1244 ? 1'h0 : T980;
  assign T980 = T1242 ? reqDoneWire_2 : T981;
  assign T981 = T1222 ? 1'h0 : T982;
  assign T982 = T1220 ? reqDoneWire_2 : T983;
  assign T983 = T1200 ? 1'h0 : T984;
  assign T984 = T1198 ? reqDoneWire_2 : T985;
  assign T985 = T1178 ? 1'h0 : T986;
  assign T986 = T1176 ? reqDoneWire_2 : T987;
  assign T987 = T1156 ? 1'h0 : T988;
  assign T988 = T1154 ? reqDoneWire_2 : T989;
  assign T989 = T1134 ? 1'h0 : T990;
  assign T990 = T1132 ? reqDoneWire_2 : T991;
  assign T991 = T1112 ? 1'h0 : T992;
  assign T992 = T1110 ? reqDoneWire_2 : T993;
  assign T993 = T1090 ? 1'h0 : T994;
  assign T994 = T1088 ? reqDoneWire_2 : T995;
  assign T995 = T1068 ? 1'h0 : T996;
  assign T996 = T1066 ? reqDoneWire_2 : T997;
  assign T997 = T86 ? 1'h0 : reqDone_2;
  assign T1003 = computeEnable & T1004;
  assign T1004 = T999 ^ 1'h1;
  assign T1005 = reqDoneWire_0 & reqDoneWire_1;
  assign reqDoneWire_1 = T1006;
  assign T1006 = T1054 ? reqDone_1 : T1007;
  assign T1007 = T1049 ? 1'h1 : T1008;
  assign T1008 = computeEnable ? reqDone_1 : 1'h0;
  assign T1049 = computeEnable & T1050;
  assign T1050 = nextRequest_1 | T1051;
  assign T1051 = ~ io_outLocValid_1;
  assign nextRequest_1 = T1052;
  assign T1052 = T1053 ? 1'h0 : io_seqProceed_1;
  assign T1053 = io_seqProceed_1 ^ 1'h1;
  assign T1675 = reset ? 1'h0 : T1009;
  assign T1009 = T1484 ? reqDoneWire_1 : T1010;
  assign T1010 = T1464 ? 1'h0 : T1011;
  assign T1011 = T1462 ? reqDoneWire_1 : T1012;
  assign T1012 = T1442 ? 1'h0 : T1013;
  assign T1013 = T1440 ? reqDoneWire_1 : T1014;
  assign T1014 = T1420 ? 1'h0 : T1015;
  assign T1015 = T1418 ? reqDoneWire_1 : T1016;
  assign T1016 = T1398 ? 1'h0 : T1017;
  assign T1017 = T1396 ? reqDoneWire_1 : T1018;
  assign T1018 = T1376 ? 1'h0 : T1019;
  assign T1019 = T1374 ? reqDoneWire_1 : T1020;
  assign T1020 = T1354 ? 1'h0 : T1021;
  assign T1021 = T1352 ? reqDoneWire_1 : T1022;
  assign T1022 = T1332 ? 1'h0 : T1023;
  assign T1023 = T1330 ? reqDoneWire_1 : T1024;
  assign T1024 = T1310 ? 1'h0 : T1025;
  assign T1025 = T1308 ? reqDoneWire_1 : T1026;
  assign T1026 = T1288 ? 1'h0 : T1027;
  assign T1027 = T1286 ? reqDoneWire_1 : T1028;
  assign T1028 = T1266 ? 1'h0 : T1029;
  assign T1029 = T1264 ? reqDoneWire_1 : T1030;
  assign T1030 = T1244 ? 1'h0 : T1031;
  assign T1031 = T1242 ? reqDoneWire_1 : T1032;
  assign T1032 = T1222 ? 1'h0 : T1033;
  assign T1033 = T1220 ? reqDoneWire_1 : T1034;
  assign T1034 = T1200 ? 1'h0 : T1035;
  assign T1035 = T1198 ? reqDoneWire_1 : T1036;
  assign T1036 = T1178 ? 1'h0 : T1037;
  assign T1037 = T1176 ? reqDoneWire_1 : T1038;
  assign T1038 = T1156 ? 1'h0 : T1039;
  assign T1039 = T1154 ? reqDoneWire_1 : T1040;
  assign T1040 = T1134 ? 1'h0 : T1041;
  assign T1041 = T1132 ? reqDoneWire_1 : T1042;
  assign T1042 = T1112 ? 1'h0 : T1043;
  assign T1043 = T1110 ? reqDoneWire_1 : T1044;
  assign T1044 = T1090 ? 1'h0 : T1045;
  assign T1045 = T1088 ? reqDoneWire_1 : T1046;
  assign T1046 = T1068 ? 1'h0 : T1047;
  assign T1047 = T1066 ? reqDoneWire_1 : T1048;
  assign T1048 = T86 ? 1'h0 : reqDone_1;
  assign T1054 = computeEnable & T1055;
  assign T1055 = T1050 ^ 1'h1;
  assign T1066 = computeEnable & T1067;
  assign T1067 = T87 ^ 1'h1;
  assign T1068 = computeEnable & T1069;
  assign T1069 = T1070 & reqDoneWire_19;
  assign T1070 = T1071 & reqDoneWire_18;
  assign T1071 = T1072 & reqDoneWire_17;
  assign T1072 = T1073 & reqDoneWire_16;
  assign T1073 = T1074 & reqDoneWire_15;
  assign T1074 = T1075 & reqDoneWire_14;
  assign T1075 = T1076 & reqDoneWire_13;
  assign T1076 = T1077 & reqDoneWire_12;
  assign T1077 = T1078 & reqDoneWire_11;
  assign T1078 = T1079 & reqDoneWire_10;
  assign T1079 = T1080 & reqDoneWire_9;
  assign T1080 = T1081 & reqDoneWire_8;
  assign T1081 = T1082 & reqDoneWire_7;
  assign T1082 = T1083 & reqDoneWire_6;
  assign T1083 = T1084 & reqDoneWire_5;
  assign T1084 = T1085 & reqDoneWire_4;
  assign T1085 = T1086 & reqDoneWire_3;
  assign T1086 = T1087 & reqDoneWire_2;
  assign T1087 = reqDoneWire_0 & reqDoneWire_1;
  assign T1088 = computeEnable & T1089;
  assign T1089 = T1069 ^ 1'h1;
  assign T1090 = computeEnable & T1091;
  assign T1091 = T1092 & reqDoneWire_19;
  assign T1092 = T1093 & reqDoneWire_18;
  assign T1093 = T1094 & reqDoneWire_17;
  assign T1094 = T1095 & reqDoneWire_16;
  assign T1095 = T1096 & reqDoneWire_15;
  assign T1096 = T1097 & reqDoneWire_14;
  assign T1097 = T1098 & reqDoneWire_13;
  assign T1098 = T1099 & reqDoneWire_12;
  assign T1099 = T1100 & reqDoneWire_11;
  assign T1100 = T1101 & reqDoneWire_10;
  assign T1101 = T1102 & reqDoneWire_9;
  assign T1102 = T1103 & reqDoneWire_8;
  assign T1103 = T1104 & reqDoneWire_7;
  assign T1104 = T1105 & reqDoneWire_6;
  assign T1105 = T1106 & reqDoneWire_5;
  assign T1106 = T1107 & reqDoneWire_4;
  assign T1107 = T1108 & reqDoneWire_3;
  assign T1108 = T1109 & reqDoneWire_2;
  assign T1109 = reqDoneWire_0 & reqDoneWire_1;
  assign T1110 = computeEnable & T1111;
  assign T1111 = T1091 ^ 1'h1;
  assign T1112 = computeEnable & T1113;
  assign T1113 = T1114 & reqDoneWire_19;
  assign T1114 = T1115 & reqDoneWire_18;
  assign T1115 = T1116 & reqDoneWire_17;
  assign T1116 = T1117 & reqDoneWire_16;
  assign T1117 = T1118 & reqDoneWire_15;
  assign T1118 = T1119 & reqDoneWire_14;
  assign T1119 = T1120 & reqDoneWire_13;
  assign T1120 = T1121 & reqDoneWire_12;
  assign T1121 = T1122 & reqDoneWire_11;
  assign T1122 = T1123 & reqDoneWire_10;
  assign T1123 = T1124 & reqDoneWire_9;
  assign T1124 = T1125 & reqDoneWire_8;
  assign T1125 = T1126 & reqDoneWire_7;
  assign T1126 = T1127 & reqDoneWire_6;
  assign T1127 = T1128 & reqDoneWire_5;
  assign T1128 = T1129 & reqDoneWire_4;
  assign T1129 = T1130 & reqDoneWire_3;
  assign T1130 = T1131 & reqDoneWire_2;
  assign T1131 = reqDoneWire_0 & reqDoneWire_1;
  assign T1132 = computeEnable & T1133;
  assign T1133 = T1113 ^ 1'h1;
  assign T1134 = computeEnable & T1135;
  assign T1135 = T1136 & reqDoneWire_19;
  assign T1136 = T1137 & reqDoneWire_18;
  assign T1137 = T1138 & reqDoneWire_17;
  assign T1138 = T1139 & reqDoneWire_16;
  assign T1139 = T1140 & reqDoneWire_15;
  assign T1140 = T1141 & reqDoneWire_14;
  assign T1141 = T1142 & reqDoneWire_13;
  assign T1142 = T1143 & reqDoneWire_12;
  assign T1143 = T1144 & reqDoneWire_11;
  assign T1144 = T1145 & reqDoneWire_10;
  assign T1145 = T1146 & reqDoneWire_9;
  assign T1146 = T1147 & reqDoneWire_8;
  assign T1147 = T1148 & reqDoneWire_7;
  assign T1148 = T1149 & reqDoneWire_6;
  assign T1149 = T1150 & reqDoneWire_5;
  assign T1150 = T1151 & reqDoneWire_4;
  assign T1151 = T1152 & reqDoneWire_3;
  assign T1152 = T1153 & reqDoneWire_2;
  assign T1153 = reqDoneWire_0 & reqDoneWire_1;
  assign T1154 = computeEnable & T1155;
  assign T1155 = T1135 ^ 1'h1;
  assign T1156 = computeEnable & T1157;
  assign T1157 = T1158 & reqDoneWire_19;
  assign T1158 = T1159 & reqDoneWire_18;
  assign T1159 = T1160 & reqDoneWire_17;
  assign T1160 = T1161 & reqDoneWire_16;
  assign T1161 = T1162 & reqDoneWire_15;
  assign T1162 = T1163 & reqDoneWire_14;
  assign T1163 = T1164 & reqDoneWire_13;
  assign T1164 = T1165 & reqDoneWire_12;
  assign T1165 = T1166 & reqDoneWire_11;
  assign T1166 = T1167 & reqDoneWire_10;
  assign T1167 = T1168 & reqDoneWire_9;
  assign T1168 = T1169 & reqDoneWire_8;
  assign T1169 = T1170 & reqDoneWire_7;
  assign T1170 = T1171 & reqDoneWire_6;
  assign T1171 = T1172 & reqDoneWire_5;
  assign T1172 = T1173 & reqDoneWire_4;
  assign T1173 = T1174 & reqDoneWire_3;
  assign T1174 = T1175 & reqDoneWire_2;
  assign T1175 = reqDoneWire_0 & reqDoneWire_1;
  assign T1176 = computeEnable & T1177;
  assign T1177 = T1157 ^ 1'h1;
  assign T1178 = computeEnable & T1179;
  assign T1179 = T1180 & reqDoneWire_19;
  assign T1180 = T1181 & reqDoneWire_18;
  assign T1181 = T1182 & reqDoneWire_17;
  assign T1182 = T1183 & reqDoneWire_16;
  assign T1183 = T1184 & reqDoneWire_15;
  assign T1184 = T1185 & reqDoneWire_14;
  assign T1185 = T1186 & reqDoneWire_13;
  assign T1186 = T1187 & reqDoneWire_12;
  assign T1187 = T1188 & reqDoneWire_11;
  assign T1188 = T1189 & reqDoneWire_10;
  assign T1189 = T1190 & reqDoneWire_9;
  assign T1190 = T1191 & reqDoneWire_8;
  assign T1191 = T1192 & reqDoneWire_7;
  assign T1192 = T1193 & reqDoneWire_6;
  assign T1193 = T1194 & reqDoneWire_5;
  assign T1194 = T1195 & reqDoneWire_4;
  assign T1195 = T1196 & reqDoneWire_3;
  assign T1196 = T1197 & reqDoneWire_2;
  assign T1197 = reqDoneWire_0 & reqDoneWire_1;
  assign T1198 = computeEnable & T1199;
  assign T1199 = T1179 ^ 1'h1;
  assign T1200 = computeEnable & T1201;
  assign T1201 = T1202 & reqDoneWire_19;
  assign T1202 = T1203 & reqDoneWire_18;
  assign T1203 = T1204 & reqDoneWire_17;
  assign T1204 = T1205 & reqDoneWire_16;
  assign T1205 = T1206 & reqDoneWire_15;
  assign T1206 = T1207 & reqDoneWire_14;
  assign T1207 = T1208 & reqDoneWire_13;
  assign T1208 = T1209 & reqDoneWire_12;
  assign T1209 = T1210 & reqDoneWire_11;
  assign T1210 = T1211 & reqDoneWire_10;
  assign T1211 = T1212 & reqDoneWire_9;
  assign T1212 = T1213 & reqDoneWire_8;
  assign T1213 = T1214 & reqDoneWire_7;
  assign T1214 = T1215 & reqDoneWire_6;
  assign T1215 = T1216 & reqDoneWire_5;
  assign T1216 = T1217 & reqDoneWire_4;
  assign T1217 = T1218 & reqDoneWire_3;
  assign T1218 = T1219 & reqDoneWire_2;
  assign T1219 = reqDoneWire_0 & reqDoneWire_1;
  assign T1220 = computeEnable & T1221;
  assign T1221 = T1201 ^ 1'h1;
  assign T1222 = computeEnable & T1223;
  assign T1223 = T1224 & reqDoneWire_19;
  assign T1224 = T1225 & reqDoneWire_18;
  assign T1225 = T1226 & reqDoneWire_17;
  assign T1226 = T1227 & reqDoneWire_16;
  assign T1227 = T1228 & reqDoneWire_15;
  assign T1228 = T1229 & reqDoneWire_14;
  assign T1229 = T1230 & reqDoneWire_13;
  assign T1230 = T1231 & reqDoneWire_12;
  assign T1231 = T1232 & reqDoneWire_11;
  assign T1232 = T1233 & reqDoneWire_10;
  assign T1233 = T1234 & reqDoneWire_9;
  assign T1234 = T1235 & reqDoneWire_8;
  assign T1235 = T1236 & reqDoneWire_7;
  assign T1236 = T1237 & reqDoneWire_6;
  assign T1237 = T1238 & reqDoneWire_5;
  assign T1238 = T1239 & reqDoneWire_4;
  assign T1239 = T1240 & reqDoneWire_3;
  assign T1240 = T1241 & reqDoneWire_2;
  assign T1241 = reqDoneWire_0 & reqDoneWire_1;
  assign T1242 = computeEnable & T1243;
  assign T1243 = T1223 ^ 1'h1;
  assign T1244 = computeEnable & T1245;
  assign T1245 = T1246 & reqDoneWire_19;
  assign T1246 = T1247 & reqDoneWire_18;
  assign T1247 = T1248 & reqDoneWire_17;
  assign T1248 = T1249 & reqDoneWire_16;
  assign T1249 = T1250 & reqDoneWire_15;
  assign T1250 = T1251 & reqDoneWire_14;
  assign T1251 = T1252 & reqDoneWire_13;
  assign T1252 = T1253 & reqDoneWire_12;
  assign T1253 = T1254 & reqDoneWire_11;
  assign T1254 = T1255 & reqDoneWire_10;
  assign T1255 = T1256 & reqDoneWire_9;
  assign T1256 = T1257 & reqDoneWire_8;
  assign T1257 = T1258 & reqDoneWire_7;
  assign T1258 = T1259 & reqDoneWire_6;
  assign T1259 = T1260 & reqDoneWire_5;
  assign T1260 = T1261 & reqDoneWire_4;
  assign T1261 = T1262 & reqDoneWire_3;
  assign T1262 = T1263 & reqDoneWire_2;
  assign T1263 = reqDoneWire_0 & reqDoneWire_1;
  assign T1264 = computeEnable & T1265;
  assign T1265 = T1245 ^ 1'h1;
  assign T1266 = computeEnable & T1267;
  assign T1267 = T1268 & reqDoneWire_19;
  assign T1268 = T1269 & reqDoneWire_18;
  assign T1269 = T1270 & reqDoneWire_17;
  assign T1270 = T1271 & reqDoneWire_16;
  assign T1271 = T1272 & reqDoneWire_15;
  assign T1272 = T1273 & reqDoneWire_14;
  assign T1273 = T1274 & reqDoneWire_13;
  assign T1274 = T1275 & reqDoneWire_12;
  assign T1275 = T1276 & reqDoneWire_11;
  assign T1276 = T1277 & reqDoneWire_10;
  assign T1277 = T1278 & reqDoneWire_9;
  assign T1278 = T1279 & reqDoneWire_8;
  assign T1279 = T1280 & reqDoneWire_7;
  assign T1280 = T1281 & reqDoneWire_6;
  assign T1281 = T1282 & reqDoneWire_5;
  assign T1282 = T1283 & reqDoneWire_4;
  assign T1283 = T1284 & reqDoneWire_3;
  assign T1284 = T1285 & reqDoneWire_2;
  assign T1285 = reqDoneWire_0 & reqDoneWire_1;
  assign T1286 = computeEnable & T1287;
  assign T1287 = T1267 ^ 1'h1;
  assign T1288 = computeEnable & T1289;
  assign T1289 = T1290 & reqDoneWire_19;
  assign T1290 = T1291 & reqDoneWire_18;
  assign T1291 = T1292 & reqDoneWire_17;
  assign T1292 = T1293 & reqDoneWire_16;
  assign T1293 = T1294 & reqDoneWire_15;
  assign T1294 = T1295 & reqDoneWire_14;
  assign T1295 = T1296 & reqDoneWire_13;
  assign T1296 = T1297 & reqDoneWire_12;
  assign T1297 = T1298 & reqDoneWire_11;
  assign T1298 = T1299 & reqDoneWire_10;
  assign T1299 = T1300 & reqDoneWire_9;
  assign T1300 = T1301 & reqDoneWire_8;
  assign T1301 = T1302 & reqDoneWire_7;
  assign T1302 = T1303 & reqDoneWire_6;
  assign T1303 = T1304 & reqDoneWire_5;
  assign T1304 = T1305 & reqDoneWire_4;
  assign T1305 = T1306 & reqDoneWire_3;
  assign T1306 = T1307 & reqDoneWire_2;
  assign T1307 = reqDoneWire_0 & reqDoneWire_1;
  assign T1308 = computeEnable & T1309;
  assign T1309 = T1289 ^ 1'h1;
  assign T1310 = computeEnable & T1311;
  assign T1311 = T1312 & reqDoneWire_19;
  assign T1312 = T1313 & reqDoneWire_18;
  assign T1313 = T1314 & reqDoneWire_17;
  assign T1314 = T1315 & reqDoneWire_16;
  assign T1315 = T1316 & reqDoneWire_15;
  assign T1316 = T1317 & reqDoneWire_14;
  assign T1317 = T1318 & reqDoneWire_13;
  assign T1318 = T1319 & reqDoneWire_12;
  assign T1319 = T1320 & reqDoneWire_11;
  assign T1320 = T1321 & reqDoneWire_10;
  assign T1321 = T1322 & reqDoneWire_9;
  assign T1322 = T1323 & reqDoneWire_8;
  assign T1323 = T1324 & reqDoneWire_7;
  assign T1324 = T1325 & reqDoneWire_6;
  assign T1325 = T1326 & reqDoneWire_5;
  assign T1326 = T1327 & reqDoneWire_4;
  assign T1327 = T1328 & reqDoneWire_3;
  assign T1328 = T1329 & reqDoneWire_2;
  assign T1329 = reqDoneWire_0 & reqDoneWire_1;
  assign T1330 = computeEnable & T1331;
  assign T1331 = T1311 ^ 1'h1;
  assign T1332 = computeEnable & T1333;
  assign T1333 = T1334 & reqDoneWire_19;
  assign T1334 = T1335 & reqDoneWire_18;
  assign T1335 = T1336 & reqDoneWire_17;
  assign T1336 = T1337 & reqDoneWire_16;
  assign T1337 = T1338 & reqDoneWire_15;
  assign T1338 = T1339 & reqDoneWire_14;
  assign T1339 = T1340 & reqDoneWire_13;
  assign T1340 = T1341 & reqDoneWire_12;
  assign T1341 = T1342 & reqDoneWire_11;
  assign T1342 = T1343 & reqDoneWire_10;
  assign T1343 = T1344 & reqDoneWire_9;
  assign T1344 = T1345 & reqDoneWire_8;
  assign T1345 = T1346 & reqDoneWire_7;
  assign T1346 = T1347 & reqDoneWire_6;
  assign T1347 = T1348 & reqDoneWire_5;
  assign T1348 = T1349 & reqDoneWire_4;
  assign T1349 = T1350 & reqDoneWire_3;
  assign T1350 = T1351 & reqDoneWire_2;
  assign T1351 = reqDoneWire_0 & reqDoneWire_1;
  assign T1352 = computeEnable & T1353;
  assign T1353 = T1333 ^ 1'h1;
  assign T1354 = computeEnable & T1355;
  assign T1355 = T1356 & reqDoneWire_19;
  assign T1356 = T1357 & reqDoneWire_18;
  assign T1357 = T1358 & reqDoneWire_17;
  assign T1358 = T1359 & reqDoneWire_16;
  assign T1359 = T1360 & reqDoneWire_15;
  assign T1360 = T1361 & reqDoneWire_14;
  assign T1361 = T1362 & reqDoneWire_13;
  assign T1362 = T1363 & reqDoneWire_12;
  assign T1363 = T1364 & reqDoneWire_11;
  assign T1364 = T1365 & reqDoneWire_10;
  assign T1365 = T1366 & reqDoneWire_9;
  assign T1366 = T1367 & reqDoneWire_8;
  assign T1367 = T1368 & reqDoneWire_7;
  assign T1368 = T1369 & reqDoneWire_6;
  assign T1369 = T1370 & reqDoneWire_5;
  assign T1370 = T1371 & reqDoneWire_4;
  assign T1371 = T1372 & reqDoneWire_3;
  assign T1372 = T1373 & reqDoneWire_2;
  assign T1373 = reqDoneWire_0 & reqDoneWire_1;
  assign T1374 = computeEnable & T1375;
  assign T1375 = T1355 ^ 1'h1;
  assign T1376 = computeEnable & T1377;
  assign T1377 = T1378 & reqDoneWire_19;
  assign T1378 = T1379 & reqDoneWire_18;
  assign T1379 = T1380 & reqDoneWire_17;
  assign T1380 = T1381 & reqDoneWire_16;
  assign T1381 = T1382 & reqDoneWire_15;
  assign T1382 = T1383 & reqDoneWire_14;
  assign T1383 = T1384 & reqDoneWire_13;
  assign T1384 = T1385 & reqDoneWire_12;
  assign T1385 = T1386 & reqDoneWire_11;
  assign T1386 = T1387 & reqDoneWire_10;
  assign T1387 = T1388 & reqDoneWire_9;
  assign T1388 = T1389 & reqDoneWire_8;
  assign T1389 = T1390 & reqDoneWire_7;
  assign T1390 = T1391 & reqDoneWire_6;
  assign T1391 = T1392 & reqDoneWire_5;
  assign T1392 = T1393 & reqDoneWire_4;
  assign T1393 = T1394 & reqDoneWire_3;
  assign T1394 = T1395 & reqDoneWire_2;
  assign T1395 = reqDoneWire_0 & reqDoneWire_1;
  assign T1396 = computeEnable & T1397;
  assign T1397 = T1377 ^ 1'h1;
  assign T1398 = computeEnable & T1399;
  assign T1399 = T1400 & reqDoneWire_19;
  assign T1400 = T1401 & reqDoneWire_18;
  assign T1401 = T1402 & reqDoneWire_17;
  assign T1402 = T1403 & reqDoneWire_16;
  assign T1403 = T1404 & reqDoneWire_15;
  assign T1404 = T1405 & reqDoneWire_14;
  assign T1405 = T1406 & reqDoneWire_13;
  assign T1406 = T1407 & reqDoneWire_12;
  assign T1407 = T1408 & reqDoneWire_11;
  assign T1408 = T1409 & reqDoneWire_10;
  assign T1409 = T1410 & reqDoneWire_9;
  assign T1410 = T1411 & reqDoneWire_8;
  assign T1411 = T1412 & reqDoneWire_7;
  assign T1412 = T1413 & reqDoneWire_6;
  assign T1413 = T1414 & reqDoneWire_5;
  assign T1414 = T1415 & reqDoneWire_4;
  assign T1415 = T1416 & reqDoneWire_3;
  assign T1416 = T1417 & reqDoneWire_2;
  assign T1417 = reqDoneWire_0 & reqDoneWire_1;
  assign T1418 = computeEnable & T1419;
  assign T1419 = T1399 ^ 1'h1;
  assign T1420 = computeEnable & T1421;
  assign T1421 = T1422 & reqDoneWire_19;
  assign T1422 = T1423 & reqDoneWire_18;
  assign T1423 = T1424 & reqDoneWire_17;
  assign T1424 = T1425 & reqDoneWire_16;
  assign T1425 = T1426 & reqDoneWire_15;
  assign T1426 = T1427 & reqDoneWire_14;
  assign T1427 = T1428 & reqDoneWire_13;
  assign T1428 = T1429 & reqDoneWire_12;
  assign T1429 = T1430 & reqDoneWire_11;
  assign T1430 = T1431 & reqDoneWire_10;
  assign T1431 = T1432 & reqDoneWire_9;
  assign T1432 = T1433 & reqDoneWire_8;
  assign T1433 = T1434 & reqDoneWire_7;
  assign T1434 = T1435 & reqDoneWire_6;
  assign T1435 = T1436 & reqDoneWire_5;
  assign T1436 = T1437 & reqDoneWire_4;
  assign T1437 = T1438 & reqDoneWire_3;
  assign T1438 = T1439 & reqDoneWire_2;
  assign T1439 = reqDoneWire_0 & reqDoneWire_1;
  assign T1440 = computeEnable & T1441;
  assign T1441 = T1421 ^ 1'h1;
  assign T1442 = computeEnable & T1443;
  assign T1443 = T1444 & reqDoneWire_19;
  assign T1444 = T1445 & reqDoneWire_18;
  assign T1445 = T1446 & reqDoneWire_17;
  assign T1446 = T1447 & reqDoneWire_16;
  assign T1447 = T1448 & reqDoneWire_15;
  assign T1448 = T1449 & reqDoneWire_14;
  assign T1449 = T1450 & reqDoneWire_13;
  assign T1450 = T1451 & reqDoneWire_12;
  assign T1451 = T1452 & reqDoneWire_11;
  assign T1452 = T1453 & reqDoneWire_10;
  assign T1453 = T1454 & reqDoneWire_9;
  assign T1454 = T1455 & reqDoneWire_8;
  assign T1455 = T1456 & reqDoneWire_7;
  assign T1456 = T1457 & reqDoneWire_6;
  assign T1457 = T1458 & reqDoneWire_5;
  assign T1458 = T1459 & reqDoneWire_4;
  assign T1459 = T1460 & reqDoneWire_3;
  assign T1460 = T1461 & reqDoneWire_2;
  assign T1461 = reqDoneWire_0 & reqDoneWire_1;
  assign T1462 = computeEnable & T1463;
  assign T1463 = T1443 ^ 1'h1;
  assign T1464 = computeEnable & T1465;
  assign T1465 = T1466 & reqDoneWire_19;
  assign T1466 = T1467 & reqDoneWire_18;
  assign T1467 = T1468 & reqDoneWire_17;
  assign T1468 = T1469 & reqDoneWire_16;
  assign T1469 = T1470 & reqDoneWire_15;
  assign T1470 = T1471 & reqDoneWire_14;
  assign T1471 = T1472 & reqDoneWire_13;
  assign T1472 = T1473 & reqDoneWire_12;
  assign T1473 = T1474 & reqDoneWire_11;
  assign T1474 = T1475 & reqDoneWire_10;
  assign T1475 = T1476 & reqDoneWire_9;
  assign T1476 = T1477 & reqDoneWire_8;
  assign T1477 = T1478 & reqDoneWire_7;
  assign T1478 = T1479 & reqDoneWire_6;
  assign T1479 = T1480 & reqDoneWire_5;
  assign T1480 = T1481 & reqDoneWire_4;
  assign T1481 = T1482 & reqDoneWire_3;
  assign T1482 = T1483 & reqDoneWire_2;
  assign T1483 = reqDoneWire_0 & reqDoneWire_1;
  assign reqDoneWire_0 = T1056;
  assign T1056 = T1064 ? reqDone_0 : T1057;
  assign T1057 = T1059 ? 1'h1 : T1058;
  assign T1058 = computeEnable ? reqDone_0 : 1'h0;
  assign T1059 = computeEnable & T1060;
  assign T1060 = nextRequest_0 | T1061;
  assign T1061 = ~ io_outLocValid_0;
  assign nextRequest_0 = T1062;
  assign T1062 = T1063 ? 1'h0 : io_seqProceed_0;
  assign T1063 = io_seqProceed_0 ^ 1'h1;
  assign T1064 = computeEnable & T1065;
  assign T1065 = T1060 ^ 1'h1;
  assign T1484 = computeEnable & T1485;
  assign T1485 = T1465 ^ 1'h1;
  assign io_seqMemAddrValid_1 = T1486;
  assign T1486 = T1487 ? 1'h1 : 1'h0;
  assign T1487 = T1488 & computeEnable;
  assign T1488 = ~ reqDone_1;
  assign io_seqMemAddrValid_2 = T1489;
  assign T1489 = T1490 ? 1'h1 : 1'h0;
  assign T1490 = T1491 & computeEnable;
  assign T1491 = ~ reqDone_2;
  assign io_seqMemAddrValid_3 = T1492;
  assign T1492 = T1493 ? 1'h1 : 1'h0;
  assign T1493 = T1494 & computeEnable;
  assign T1494 = ~ reqDone_3;
  assign io_seqMemAddrValid_4 = T1495;
  assign T1495 = T1496 ? 1'h1 : 1'h0;
  assign T1496 = T1497 & computeEnable;
  assign T1497 = ~ reqDone_4;
  assign io_seqMemAddrValid_5 = T1498;
  assign T1498 = T1499 ? 1'h1 : 1'h0;
  assign T1499 = T1500 & computeEnable;
  assign T1500 = ~ reqDone_5;
  assign io_seqMemAddrValid_6 = T1501;
  assign T1501 = T1502 ? 1'h1 : 1'h0;
  assign T1502 = T1503 & computeEnable;
  assign T1503 = ~ reqDone_6;
  assign io_seqMemAddrValid_7 = T1504;
  assign T1504 = T1505 ? 1'h1 : 1'h0;
  assign T1505 = T1506 & computeEnable;
  assign T1506 = ~ reqDone_7;
  assign io_seqMemAddrValid_8 = T1507;
  assign T1507 = T1508 ? 1'h1 : 1'h0;
  assign T1508 = T1509 & computeEnable;
  assign T1509 = ~ reqDone_8;
  assign io_seqMemAddrValid_9 = T1510;
  assign T1510 = T1511 ? 1'h1 : 1'h0;
  assign T1511 = T1512 & computeEnable;
  assign T1512 = ~ reqDone_9;
  assign io_seqMemAddrValid_10 = T1513;
  assign T1513 = T1514 ? 1'h1 : 1'h0;
  assign T1514 = T1515 & computeEnable;
  assign T1515 = ~ reqDone_10;
  assign io_seqMemAddrValid_11 = T1516;
  assign T1516 = T1517 ? 1'h1 : 1'h0;
  assign T1517 = T1518 & computeEnable;
  assign T1518 = ~ reqDone_11;
  assign io_seqMemAddrValid_12 = T1519;
  assign T1519 = T1520 ? 1'h1 : 1'h0;
  assign T1520 = T1521 & computeEnable;
  assign T1521 = ~ reqDone_12;
  assign io_seqMemAddrValid_13 = T1522;
  assign T1522 = T1523 ? 1'h1 : 1'h0;
  assign T1523 = T1524 & computeEnable;
  assign T1524 = ~ reqDone_13;
  assign io_seqMemAddrValid_14 = T1525;
  assign T1525 = T1526 ? 1'h1 : 1'h0;
  assign T1526 = T1527 & computeEnable;
  assign T1527 = ~ reqDone_14;
  assign io_seqMemAddrValid_15 = T1528;
  assign T1528 = T1529 ? 1'h1 : 1'h0;
  assign T1529 = T1530 & computeEnable;
  assign T1530 = ~ reqDone_15;
  assign io_seqMemAddrValid_16 = T1531;
  assign T1531 = T1532 ? 1'h1 : 1'h0;
  assign T1532 = T1533 & computeEnable;
  assign T1533 = ~ reqDone_16;
  assign io_seqMemAddrValid_17 = T1534;
  assign T1534 = T1535 ? 1'h1 : 1'h0;
  assign T1535 = T1536 & computeEnable;
  assign T1536 = ~ reqDone_17;
  assign io_seqMemAddrValid_18 = T1537;
  assign T1537 = T1538 ? 1'h1 : 1'h0;
  assign T1538 = T1539 & computeEnable;
  assign T1539 = ~ reqDone_18;
  assign io_seqMemAddrValid_19 = T1540;
  assign T1540 = T1541 ? 1'h1 : 1'h0;
  assign T1541 = T1542 & computeEnable;
  assign T1542 = ~ reqDone_19;
  assign io_seqMemAddr_0 = T1543;
  assign T1543 = T1 ? seqMemAddr : seqMemAddr;
  assign T1676 = T1677[4'h8:1'h0];
  assign T1677 = reset ? 514'h0 : T1544;
  assign T1544 = T1623 ? T1687 : T1545;
  assign T1545 = T1615 ? ssEnd : T1678;
  assign T1678 = {505'h0, T1546};
  assign T1546 = T1613 ? T1612 : T1547;
  assign T1547 = T1590 ? prologueDepth : T1548;
  assign T1548 = T1549 ? 9'h0 : seqMemAddr;
  assign T1549 = T1550 & startComputeValid;
  assign T1550 = startComputeValid | nextSeqRdy;
  assign nextSeqRdy = T1551;
  assign T1551 = T1484 ? 1'h0 : T1552;
  assign T1552 = T1464 ? 1'h1 : T1553;
  assign T1553 = T1462 ? 1'h0 : T1554;
  assign T1554 = T1442 ? 1'h1 : T1555;
  assign T1555 = T1440 ? 1'h0 : T1556;
  assign T1556 = T1420 ? 1'h1 : T1557;
  assign T1557 = T1418 ? 1'h0 : T1558;
  assign T1558 = T1398 ? 1'h1 : T1559;
  assign T1559 = T1396 ? 1'h0 : T1560;
  assign T1560 = T1376 ? 1'h1 : T1561;
  assign T1561 = T1374 ? 1'h0 : T1562;
  assign T1562 = T1354 ? 1'h1 : T1563;
  assign T1563 = T1352 ? 1'h0 : T1564;
  assign T1564 = T1332 ? 1'h1 : T1565;
  assign T1565 = T1330 ? 1'h0 : T1566;
  assign T1566 = T1310 ? 1'h1 : T1567;
  assign T1567 = T1308 ? 1'h0 : T1568;
  assign T1568 = T1288 ? 1'h1 : T1569;
  assign T1569 = T1286 ? 1'h0 : T1570;
  assign T1570 = T1266 ? 1'h1 : T1571;
  assign T1571 = T1264 ? 1'h0 : T1572;
  assign T1572 = T1244 ? 1'h1 : T1573;
  assign T1573 = T1242 ? 1'h0 : T1574;
  assign T1574 = T1222 ? 1'h1 : T1575;
  assign T1575 = T1220 ? 1'h0 : T1576;
  assign T1576 = T1200 ? 1'h1 : T1577;
  assign T1577 = T1198 ? 1'h0 : T1578;
  assign T1578 = T1178 ? 1'h1 : T1579;
  assign T1579 = T1176 ? 1'h0 : T1580;
  assign T1580 = T1156 ? 1'h1 : T1581;
  assign T1581 = T1154 ? 1'h0 : T1582;
  assign T1582 = T1134 ? 1'h1 : T1583;
  assign T1583 = T1132 ? 1'h0 : T1584;
  assign T1584 = T1112 ? 1'h1 : T1585;
  assign T1585 = T1110 ? 1'h0 : T1586;
  assign T1586 = T1090 ? 1'h1 : T1587;
  assign T1587 = T1088 ? 1'h0 : T1588;
  assign T1588 = T1068 ? 1'h1 : T1589;
  assign T1589 = T1066 ? 1'h0 : T86;
  assign T1590 = T1607 & T1591;
  assign T1591 = T1595 | T1592;
  assign T1592 = epilogueSpill != 9'h0;
  assign T1679 = T1680[4'h8:1'h0];
  assign T1680 = reset ? 10'h0 : T1593;
  assign T1593 = T11 ? T1594 : T1681;
  assign T1681 = {1'h0, epilogueSpill};
  assign T1594 = io_inConfig[5'h10:3'h7];
  assign T1595 = currentIter < T1596;
  assign T1596 = iterCount - 32'h1;
  assign T1682 = reset ? 32'h0 : T1597;
  assign T1597 = T1599 ? T1683 : iterCount;
  assign T1683 = {13'h0, T1598};
  assign T1598 = io_inConfig[5'h12:1'h0];
  assign T1599 = T21 & T1600;
  assign T1600 = T1603 & T1601;
  assign T1601 = T1602 == 3'h1;
  assign T1602 = io_inConfig[5'h15:5'h13];
  assign T1603 = T19 ^ 1'h1;
  assign T1684 = reset ? 32'h0 : T1604;
  assign T1604 = T1590 ? T1606 : T1605;
  assign T1605 = T1549 ? 32'h0 : currentIter;
  assign T1606 = currentIter + 32'h1;
  assign T1607 = T1610 & T1608;
  assign T1608 = T1685 == T1609;
  assign T1609 = ssEnd - 514'h1;
  assign T1685 = {505'h0, seqMemAddr};
  assign T1610 = T1550 & T1611;
  assign T1611 = startComputeValid ^ 1'h1;
  assign T1612 = seqMemAddr + 9'h1;
  assign T1613 = T1607 & T1614;
  assign T1614 = T1591 ^ 1'h1;
  assign T1615 = T1610 & T1616;
  assign T1616 = T1621 & T1617;
  assign T1617 = T1620 & T1618;
  assign T1618 = T1686 == T1619;
  assign T1619 = ssEnd - 514'h1;
  assign T1686 = {505'h0, seqMemAddr};
  assign T1620 = currentIter == iterCount;
  assign T1621 = T1608 ^ 1'h1;
  assign T1687 = {505'h0, T1622};
  assign T1622 = seqMemAddr + 9'h1;
  assign T1623 = T1610 & T1624;
  assign T1624 = T1625 ^ 1'h1;
  assign T1625 = T1608 | T1617;
  assign io_seqMemAddr_1 = T1626;
  assign T1626 = T1487 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_2 = T1627;
  assign T1627 = T1490 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_3 = T1628;
  assign T1628 = T1493 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_4 = T1629;
  assign T1629 = T1496 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_5 = T1630;
  assign T1630 = T1499 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_6 = T1631;
  assign T1631 = T1502 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_7 = T1632;
  assign T1632 = T1505 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_8 = T1633;
  assign T1633 = T1508 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_9 = T1634;
  assign T1634 = T1511 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_10 = T1635;
  assign T1635 = T1514 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_11 = T1636;
  assign T1636 = T1517 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_12 = T1637;
  assign T1637 = T1520 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_13 = T1638;
  assign T1638 = T1523 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_14 = T1639;
  assign T1639 = T1526 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_15 = T1640;
  assign T1640 = T1529 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_16 = T1641;
  assign T1641 = T1532 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_17 = T1642;
  assign T1642 = T1535 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_18 = T1643;
  assign T1643 = T1538 ? seqMemAddr : seqMemAddr;
  assign io_seqMemAddr_19 = T1644;
  assign T1644 = T1541 ? seqMemAddr : seqMemAddr;
  controllerConfigure_0 fabOutSeqCtrlConfigure(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       //.io_outConfig(  )
       //.io_outValid(  )
       .io_computeCtrl( fabOutSeqCtrlConfigure_io_computeCtrl ),
       .io_computeCtrlValid( fabOutSeqCtrlConfigure_io_computeCtrlValid )
  );

  always @(posedge clk) begin
    if(reset) begin
      computeEnable <= 1'h0;
    end else if(T42) begin
      computeEnable <= 1'h0;
    end else if(T39) begin
      computeEnable <= 1'h0;
    end else if(T5) begin
      computeEnable <= 1'h1;
    end
    if(reset) begin
      epilogueDepth <= 9'h0;
    end else if(T11) begin
      epilogueDepth <= T1649;
    end
    steadyStateDepth <= T1651;
    if(reset) begin
      prologueDepth <= 9'h0;
    end else if(T27) begin
      prologueDepth <= T1655;
    end
    if(reset) begin
      reqDone_0 <= 1'h0;
    end else if(T1484) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1464) begin
      reqDone_0 <= 1'h0;
    end else if(T1462) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1442) begin
      reqDone_0 <= 1'h0;
    end else if(T1440) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1420) begin
      reqDone_0 <= 1'h0;
    end else if(T1418) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1398) begin
      reqDone_0 <= 1'h0;
    end else if(T1396) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1376) begin
      reqDone_0 <= 1'h0;
    end else if(T1374) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1354) begin
      reqDone_0 <= 1'h0;
    end else if(T1352) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1332) begin
      reqDone_0 <= 1'h0;
    end else if(T1330) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1310) begin
      reqDone_0 <= 1'h0;
    end else if(T1308) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1288) begin
      reqDone_0 <= 1'h0;
    end else if(T1286) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1266) begin
      reqDone_0 <= 1'h0;
    end else if(T1264) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1244) begin
      reqDone_0 <= 1'h0;
    end else if(T1242) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1222) begin
      reqDone_0 <= 1'h0;
    end else if(T1220) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1200) begin
      reqDone_0 <= 1'h0;
    end else if(T1198) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1178) begin
      reqDone_0 <= 1'h0;
    end else if(T1176) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1156) begin
      reqDone_0 <= 1'h0;
    end else if(T1154) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1134) begin
      reqDone_0 <= 1'h0;
    end else if(T1132) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1112) begin
      reqDone_0 <= 1'h0;
    end else if(T1110) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1090) begin
      reqDone_0 <= 1'h0;
    end else if(T1088) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T1068) begin
      reqDone_0 <= 1'h0;
    end else if(T1066) begin
      reqDone_0 <= reqDoneWire_0;
    end else if(T86) begin
      reqDone_0 <= 1'h0;
    end
    if(reset) begin
      reqDone_19 <= 1'h0;
    end else if(T1484) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1464) begin
      reqDone_19 <= 1'h0;
    end else if(T1462) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1442) begin
      reqDone_19 <= 1'h0;
    end else if(T1440) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1420) begin
      reqDone_19 <= 1'h0;
    end else if(T1418) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1398) begin
      reqDone_19 <= 1'h0;
    end else if(T1396) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1376) begin
      reqDone_19 <= 1'h0;
    end else if(T1374) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1354) begin
      reqDone_19 <= 1'h0;
    end else if(T1352) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1332) begin
      reqDone_19 <= 1'h0;
    end else if(T1330) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1310) begin
      reqDone_19 <= 1'h0;
    end else if(T1308) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1288) begin
      reqDone_19 <= 1'h0;
    end else if(T1286) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1266) begin
      reqDone_19 <= 1'h0;
    end else if(T1264) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1244) begin
      reqDone_19 <= 1'h0;
    end else if(T1242) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1222) begin
      reqDone_19 <= 1'h0;
    end else if(T1220) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1200) begin
      reqDone_19 <= 1'h0;
    end else if(T1198) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1178) begin
      reqDone_19 <= 1'h0;
    end else if(T1176) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1156) begin
      reqDone_19 <= 1'h0;
    end else if(T1154) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1134) begin
      reqDone_19 <= 1'h0;
    end else if(T1132) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1112) begin
      reqDone_19 <= 1'h0;
    end else if(T1110) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1090) begin
      reqDone_19 <= 1'h0;
    end else if(T1088) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T1068) begin
      reqDone_19 <= 1'h0;
    end else if(T1066) begin
      reqDone_19 <= reqDoneWire_19;
    end else if(T86) begin
      reqDone_19 <= 1'h0;
    end
    if(reset) begin
      reqDone_18 <= 1'h0;
    end else if(T1484) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1464) begin
      reqDone_18 <= 1'h0;
    end else if(T1462) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1442) begin
      reqDone_18 <= 1'h0;
    end else if(T1440) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1420) begin
      reqDone_18 <= 1'h0;
    end else if(T1418) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1398) begin
      reqDone_18 <= 1'h0;
    end else if(T1396) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1376) begin
      reqDone_18 <= 1'h0;
    end else if(T1374) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1354) begin
      reqDone_18 <= 1'h0;
    end else if(T1352) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1332) begin
      reqDone_18 <= 1'h0;
    end else if(T1330) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1310) begin
      reqDone_18 <= 1'h0;
    end else if(T1308) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1288) begin
      reqDone_18 <= 1'h0;
    end else if(T1286) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1266) begin
      reqDone_18 <= 1'h0;
    end else if(T1264) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1244) begin
      reqDone_18 <= 1'h0;
    end else if(T1242) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1222) begin
      reqDone_18 <= 1'h0;
    end else if(T1220) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1200) begin
      reqDone_18 <= 1'h0;
    end else if(T1198) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1178) begin
      reqDone_18 <= 1'h0;
    end else if(T1176) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1156) begin
      reqDone_18 <= 1'h0;
    end else if(T1154) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1134) begin
      reqDone_18 <= 1'h0;
    end else if(T1132) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1112) begin
      reqDone_18 <= 1'h0;
    end else if(T1110) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1090) begin
      reqDone_18 <= 1'h0;
    end else if(T1088) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T1068) begin
      reqDone_18 <= 1'h0;
    end else if(T1066) begin
      reqDone_18 <= reqDoneWire_18;
    end else if(T86) begin
      reqDone_18 <= 1'h0;
    end
    if(reset) begin
      reqDone_17 <= 1'h0;
    end else if(T1484) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1464) begin
      reqDone_17 <= 1'h0;
    end else if(T1462) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1442) begin
      reqDone_17 <= 1'h0;
    end else if(T1440) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1420) begin
      reqDone_17 <= 1'h0;
    end else if(T1418) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1398) begin
      reqDone_17 <= 1'h0;
    end else if(T1396) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1376) begin
      reqDone_17 <= 1'h0;
    end else if(T1374) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1354) begin
      reqDone_17 <= 1'h0;
    end else if(T1352) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1332) begin
      reqDone_17 <= 1'h0;
    end else if(T1330) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1310) begin
      reqDone_17 <= 1'h0;
    end else if(T1308) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1288) begin
      reqDone_17 <= 1'h0;
    end else if(T1286) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1266) begin
      reqDone_17 <= 1'h0;
    end else if(T1264) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1244) begin
      reqDone_17 <= 1'h0;
    end else if(T1242) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1222) begin
      reqDone_17 <= 1'h0;
    end else if(T1220) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1200) begin
      reqDone_17 <= 1'h0;
    end else if(T1198) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1178) begin
      reqDone_17 <= 1'h0;
    end else if(T1176) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1156) begin
      reqDone_17 <= 1'h0;
    end else if(T1154) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1134) begin
      reqDone_17 <= 1'h0;
    end else if(T1132) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1112) begin
      reqDone_17 <= 1'h0;
    end else if(T1110) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1090) begin
      reqDone_17 <= 1'h0;
    end else if(T1088) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T1068) begin
      reqDone_17 <= 1'h0;
    end else if(T1066) begin
      reqDone_17 <= reqDoneWire_17;
    end else if(T86) begin
      reqDone_17 <= 1'h0;
    end
    if(reset) begin
      reqDone_16 <= 1'h0;
    end else if(T1484) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1464) begin
      reqDone_16 <= 1'h0;
    end else if(T1462) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1442) begin
      reqDone_16 <= 1'h0;
    end else if(T1440) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1420) begin
      reqDone_16 <= 1'h0;
    end else if(T1418) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1398) begin
      reqDone_16 <= 1'h0;
    end else if(T1396) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1376) begin
      reqDone_16 <= 1'h0;
    end else if(T1374) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1354) begin
      reqDone_16 <= 1'h0;
    end else if(T1352) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1332) begin
      reqDone_16 <= 1'h0;
    end else if(T1330) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1310) begin
      reqDone_16 <= 1'h0;
    end else if(T1308) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1288) begin
      reqDone_16 <= 1'h0;
    end else if(T1286) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1266) begin
      reqDone_16 <= 1'h0;
    end else if(T1264) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1244) begin
      reqDone_16 <= 1'h0;
    end else if(T1242) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1222) begin
      reqDone_16 <= 1'h0;
    end else if(T1220) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1200) begin
      reqDone_16 <= 1'h0;
    end else if(T1198) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1178) begin
      reqDone_16 <= 1'h0;
    end else if(T1176) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1156) begin
      reqDone_16 <= 1'h0;
    end else if(T1154) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1134) begin
      reqDone_16 <= 1'h0;
    end else if(T1132) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1112) begin
      reqDone_16 <= 1'h0;
    end else if(T1110) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1090) begin
      reqDone_16 <= 1'h0;
    end else if(T1088) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T1068) begin
      reqDone_16 <= 1'h0;
    end else if(T1066) begin
      reqDone_16 <= reqDoneWire_16;
    end else if(T86) begin
      reqDone_16 <= 1'h0;
    end
    if(reset) begin
      reqDone_15 <= 1'h0;
    end else if(T1484) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1464) begin
      reqDone_15 <= 1'h0;
    end else if(T1462) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1442) begin
      reqDone_15 <= 1'h0;
    end else if(T1440) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1420) begin
      reqDone_15 <= 1'h0;
    end else if(T1418) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1398) begin
      reqDone_15 <= 1'h0;
    end else if(T1396) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1376) begin
      reqDone_15 <= 1'h0;
    end else if(T1374) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1354) begin
      reqDone_15 <= 1'h0;
    end else if(T1352) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1332) begin
      reqDone_15 <= 1'h0;
    end else if(T1330) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1310) begin
      reqDone_15 <= 1'h0;
    end else if(T1308) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1288) begin
      reqDone_15 <= 1'h0;
    end else if(T1286) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1266) begin
      reqDone_15 <= 1'h0;
    end else if(T1264) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1244) begin
      reqDone_15 <= 1'h0;
    end else if(T1242) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1222) begin
      reqDone_15 <= 1'h0;
    end else if(T1220) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1200) begin
      reqDone_15 <= 1'h0;
    end else if(T1198) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1178) begin
      reqDone_15 <= 1'h0;
    end else if(T1176) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1156) begin
      reqDone_15 <= 1'h0;
    end else if(T1154) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1134) begin
      reqDone_15 <= 1'h0;
    end else if(T1132) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1112) begin
      reqDone_15 <= 1'h0;
    end else if(T1110) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1090) begin
      reqDone_15 <= 1'h0;
    end else if(T1088) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T1068) begin
      reqDone_15 <= 1'h0;
    end else if(T1066) begin
      reqDone_15 <= reqDoneWire_15;
    end else if(T86) begin
      reqDone_15 <= 1'h0;
    end
    if(reset) begin
      reqDone_14 <= 1'h0;
    end else if(T1484) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1464) begin
      reqDone_14 <= 1'h0;
    end else if(T1462) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1442) begin
      reqDone_14 <= 1'h0;
    end else if(T1440) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1420) begin
      reqDone_14 <= 1'h0;
    end else if(T1418) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1398) begin
      reqDone_14 <= 1'h0;
    end else if(T1396) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1376) begin
      reqDone_14 <= 1'h0;
    end else if(T1374) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1354) begin
      reqDone_14 <= 1'h0;
    end else if(T1352) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1332) begin
      reqDone_14 <= 1'h0;
    end else if(T1330) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1310) begin
      reqDone_14 <= 1'h0;
    end else if(T1308) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1288) begin
      reqDone_14 <= 1'h0;
    end else if(T1286) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1266) begin
      reqDone_14 <= 1'h0;
    end else if(T1264) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1244) begin
      reqDone_14 <= 1'h0;
    end else if(T1242) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1222) begin
      reqDone_14 <= 1'h0;
    end else if(T1220) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1200) begin
      reqDone_14 <= 1'h0;
    end else if(T1198) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1178) begin
      reqDone_14 <= 1'h0;
    end else if(T1176) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1156) begin
      reqDone_14 <= 1'h0;
    end else if(T1154) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1134) begin
      reqDone_14 <= 1'h0;
    end else if(T1132) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1112) begin
      reqDone_14 <= 1'h0;
    end else if(T1110) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1090) begin
      reqDone_14 <= 1'h0;
    end else if(T1088) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T1068) begin
      reqDone_14 <= 1'h0;
    end else if(T1066) begin
      reqDone_14 <= reqDoneWire_14;
    end else if(T86) begin
      reqDone_14 <= 1'h0;
    end
    if(reset) begin
      reqDone_13 <= 1'h0;
    end else if(T1484) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1464) begin
      reqDone_13 <= 1'h0;
    end else if(T1462) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1442) begin
      reqDone_13 <= 1'h0;
    end else if(T1440) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1420) begin
      reqDone_13 <= 1'h0;
    end else if(T1418) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1398) begin
      reqDone_13 <= 1'h0;
    end else if(T1396) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1376) begin
      reqDone_13 <= 1'h0;
    end else if(T1374) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1354) begin
      reqDone_13 <= 1'h0;
    end else if(T1352) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1332) begin
      reqDone_13 <= 1'h0;
    end else if(T1330) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1310) begin
      reqDone_13 <= 1'h0;
    end else if(T1308) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1288) begin
      reqDone_13 <= 1'h0;
    end else if(T1286) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1266) begin
      reqDone_13 <= 1'h0;
    end else if(T1264) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1244) begin
      reqDone_13 <= 1'h0;
    end else if(T1242) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1222) begin
      reqDone_13 <= 1'h0;
    end else if(T1220) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1200) begin
      reqDone_13 <= 1'h0;
    end else if(T1198) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1178) begin
      reqDone_13 <= 1'h0;
    end else if(T1176) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1156) begin
      reqDone_13 <= 1'h0;
    end else if(T1154) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1134) begin
      reqDone_13 <= 1'h0;
    end else if(T1132) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1112) begin
      reqDone_13 <= 1'h0;
    end else if(T1110) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1090) begin
      reqDone_13 <= 1'h0;
    end else if(T1088) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T1068) begin
      reqDone_13 <= 1'h0;
    end else if(T1066) begin
      reqDone_13 <= reqDoneWire_13;
    end else if(T86) begin
      reqDone_13 <= 1'h0;
    end
    if(reset) begin
      reqDone_12 <= 1'h0;
    end else if(T1484) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1464) begin
      reqDone_12 <= 1'h0;
    end else if(T1462) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1442) begin
      reqDone_12 <= 1'h0;
    end else if(T1440) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1420) begin
      reqDone_12 <= 1'h0;
    end else if(T1418) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1398) begin
      reqDone_12 <= 1'h0;
    end else if(T1396) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1376) begin
      reqDone_12 <= 1'h0;
    end else if(T1374) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1354) begin
      reqDone_12 <= 1'h0;
    end else if(T1352) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1332) begin
      reqDone_12 <= 1'h0;
    end else if(T1330) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1310) begin
      reqDone_12 <= 1'h0;
    end else if(T1308) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1288) begin
      reqDone_12 <= 1'h0;
    end else if(T1286) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1266) begin
      reqDone_12 <= 1'h0;
    end else if(T1264) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1244) begin
      reqDone_12 <= 1'h0;
    end else if(T1242) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1222) begin
      reqDone_12 <= 1'h0;
    end else if(T1220) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1200) begin
      reqDone_12 <= 1'h0;
    end else if(T1198) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1178) begin
      reqDone_12 <= 1'h0;
    end else if(T1176) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1156) begin
      reqDone_12 <= 1'h0;
    end else if(T1154) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1134) begin
      reqDone_12 <= 1'h0;
    end else if(T1132) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1112) begin
      reqDone_12 <= 1'h0;
    end else if(T1110) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1090) begin
      reqDone_12 <= 1'h0;
    end else if(T1088) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T1068) begin
      reqDone_12 <= 1'h0;
    end else if(T1066) begin
      reqDone_12 <= reqDoneWire_12;
    end else if(T86) begin
      reqDone_12 <= 1'h0;
    end
    if(reset) begin
      reqDone_11 <= 1'h0;
    end else if(T1484) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1464) begin
      reqDone_11 <= 1'h0;
    end else if(T1462) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1442) begin
      reqDone_11 <= 1'h0;
    end else if(T1440) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1420) begin
      reqDone_11 <= 1'h0;
    end else if(T1418) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1398) begin
      reqDone_11 <= 1'h0;
    end else if(T1396) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1376) begin
      reqDone_11 <= 1'h0;
    end else if(T1374) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1354) begin
      reqDone_11 <= 1'h0;
    end else if(T1352) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1332) begin
      reqDone_11 <= 1'h0;
    end else if(T1330) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1310) begin
      reqDone_11 <= 1'h0;
    end else if(T1308) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1288) begin
      reqDone_11 <= 1'h0;
    end else if(T1286) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1266) begin
      reqDone_11 <= 1'h0;
    end else if(T1264) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1244) begin
      reqDone_11 <= 1'h0;
    end else if(T1242) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1222) begin
      reqDone_11 <= 1'h0;
    end else if(T1220) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1200) begin
      reqDone_11 <= 1'h0;
    end else if(T1198) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1178) begin
      reqDone_11 <= 1'h0;
    end else if(T1176) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1156) begin
      reqDone_11 <= 1'h0;
    end else if(T1154) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1134) begin
      reqDone_11 <= 1'h0;
    end else if(T1132) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1112) begin
      reqDone_11 <= 1'h0;
    end else if(T1110) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1090) begin
      reqDone_11 <= 1'h0;
    end else if(T1088) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T1068) begin
      reqDone_11 <= 1'h0;
    end else if(T1066) begin
      reqDone_11 <= reqDoneWire_11;
    end else if(T86) begin
      reqDone_11 <= 1'h0;
    end
    if(reset) begin
      reqDone_10 <= 1'h0;
    end else if(T1484) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1464) begin
      reqDone_10 <= 1'h0;
    end else if(T1462) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1442) begin
      reqDone_10 <= 1'h0;
    end else if(T1440) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1420) begin
      reqDone_10 <= 1'h0;
    end else if(T1418) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1398) begin
      reqDone_10 <= 1'h0;
    end else if(T1396) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1376) begin
      reqDone_10 <= 1'h0;
    end else if(T1374) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1354) begin
      reqDone_10 <= 1'h0;
    end else if(T1352) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1332) begin
      reqDone_10 <= 1'h0;
    end else if(T1330) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1310) begin
      reqDone_10 <= 1'h0;
    end else if(T1308) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1288) begin
      reqDone_10 <= 1'h0;
    end else if(T1286) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1266) begin
      reqDone_10 <= 1'h0;
    end else if(T1264) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1244) begin
      reqDone_10 <= 1'h0;
    end else if(T1242) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1222) begin
      reqDone_10 <= 1'h0;
    end else if(T1220) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1200) begin
      reqDone_10 <= 1'h0;
    end else if(T1198) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1178) begin
      reqDone_10 <= 1'h0;
    end else if(T1176) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1156) begin
      reqDone_10 <= 1'h0;
    end else if(T1154) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1134) begin
      reqDone_10 <= 1'h0;
    end else if(T1132) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1112) begin
      reqDone_10 <= 1'h0;
    end else if(T1110) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1090) begin
      reqDone_10 <= 1'h0;
    end else if(T1088) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T1068) begin
      reqDone_10 <= 1'h0;
    end else if(T1066) begin
      reqDone_10 <= reqDoneWire_10;
    end else if(T86) begin
      reqDone_10 <= 1'h0;
    end
    if(reset) begin
      reqDone_9 <= 1'h0;
    end else if(T1484) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1464) begin
      reqDone_9 <= 1'h0;
    end else if(T1462) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1442) begin
      reqDone_9 <= 1'h0;
    end else if(T1440) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1420) begin
      reqDone_9 <= 1'h0;
    end else if(T1418) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1398) begin
      reqDone_9 <= 1'h0;
    end else if(T1396) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1376) begin
      reqDone_9 <= 1'h0;
    end else if(T1374) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1354) begin
      reqDone_9 <= 1'h0;
    end else if(T1352) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1332) begin
      reqDone_9 <= 1'h0;
    end else if(T1330) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1310) begin
      reqDone_9 <= 1'h0;
    end else if(T1308) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1288) begin
      reqDone_9 <= 1'h0;
    end else if(T1286) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1266) begin
      reqDone_9 <= 1'h0;
    end else if(T1264) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1244) begin
      reqDone_9 <= 1'h0;
    end else if(T1242) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1222) begin
      reqDone_9 <= 1'h0;
    end else if(T1220) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1200) begin
      reqDone_9 <= 1'h0;
    end else if(T1198) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1178) begin
      reqDone_9 <= 1'h0;
    end else if(T1176) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1156) begin
      reqDone_9 <= 1'h0;
    end else if(T1154) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1134) begin
      reqDone_9 <= 1'h0;
    end else if(T1132) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1112) begin
      reqDone_9 <= 1'h0;
    end else if(T1110) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1090) begin
      reqDone_9 <= 1'h0;
    end else if(T1088) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T1068) begin
      reqDone_9 <= 1'h0;
    end else if(T1066) begin
      reqDone_9 <= reqDoneWire_9;
    end else if(T86) begin
      reqDone_9 <= 1'h0;
    end
    if(reset) begin
      reqDone_8 <= 1'h0;
    end else if(T1484) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1464) begin
      reqDone_8 <= 1'h0;
    end else if(T1462) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1442) begin
      reqDone_8 <= 1'h0;
    end else if(T1440) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1420) begin
      reqDone_8 <= 1'h0;
    end else if(T1418) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1398) begin
      reqDone_8 <= 1'h0;
    end else if(T1396) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1376) begin
      reqDone_8 <= 1'h0;
    end else if(T1374) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1354) begin
      reqDone_8 <= 1'h0;
    end else if(T1352) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1332) begin
      reqDone_8 <= 1'h0;
    end else if(T1330) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1310) begin
      reqDone_8 <= 1'h0;
    end else if(T1308) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1288) begin
      reqDone_8 <= 1'h0;
    end else if(T1286) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1266) begin
      reqDone_8 <= 1'h0;
    end else if(T1264) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1244) begin
      reqDone_8 <= 1'h0;
    end else if(T1242) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1222) begin
      reqDone_8 <= 1'h0;
    end else if(T1220) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1200) begin
      reqDone_8 <= 1'h0;
    end else if(T1198) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1178) begin
      reqDone_8 <= 1'h0;
    end else if(T1176) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1156) begin
      reqDone_8 <= 1'h0;
    end else if(T1154) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1134) begin
      reqDone_8 <= 1'h0;
    end else if(T1132) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1112) begin
      reqDone_8 <= 1'h0;
    end else if(T1110) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1090) begin
      reqDone_8 <= 1'h0;
    end else if(T1088) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T1068) begin
      reqDone_8 <= 1'h0;
    end else if(T1066) begin
      reqDone_8 <= reqDoneWire_8;
    end else if(T86) begin
      reqDone_8 <= 1'h0;
    end
    if(reset) begin
      reqDone_7 <= 1'h0;
    end else if(T1484) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1464) begin
      reqDone_7 <= 1'h0;
    end else if(T1462) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1442) begin
      reqDone_7 <= 1'h0;
    end else if(T1440) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1420) begin
      reqDone_7 <= 1'h0;
    end else if(T1418) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1398) begin
      reqDone_7 <= 1'h0;
    end else if(T1396) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1376) begin
      reqDone_7 <= 1'h0;
    end else if(T1374) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1354) begin
      reqDone_7 <= 1'h0;
    end else if(T1352) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1332) begin
      reqDone_7 <= 1'h0;
    end else if(T1330) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1310) begin
      reqDone_7 <= 1'h0;
    end else if(T1308) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1288) begin
      reqDone_7 <= 1'h0;
    end else if(T1286) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1266) begin
      reqDone_7 <= 1'h0;
    end else if(T1264) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1244) begin
      reqDone_7 <= 1'h0;
    end else if(T1242) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1222) begin
      reqDone_7 <= 1'h0;
    end else if(T1220) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1200) begin
      reqDone_7 <= 1'h0;
    end else if(T1198) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1178) begin
      reqDone_7 <= 1'h0;
    end else if(T1176) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1156) begin
      reqDone_7 <= 1'h0;
    end else if(T1154) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1134) begin
      reqDone_7 <= 1'h0;
    end else if(T1132) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1112) begin
      reqDone_7 <= 1'h0;
    end else if(T1110) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1090) begin
      reqDone_7 <= 1'h0;
    end else if(T1088) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T1068) begin
      reqDone_7 <= 1'h0;
    end else if(T1066) begin
      reqDone_7 <= reqDoneWire_7;
    end else if(T86) begin
      reqDone_7 <= 1'h0;
    end
    if(reset) begin
      reqDone_6 <= 1'h0;
    end else if(T1484) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1464) begin
      reqDone_6 <= 1'h0;
    end else if(T1462) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1442) begin
      reqDone_6 <= 1'h0;
    end else if(T1440) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1420) begin
      reqDone_6 <= 1'h0;
    end else if(T1418) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1398) begin
      reqDone_6 <= 1'h0;
    end else if(T1396) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1376) begin
      reqDone_6 <= 1'h0;
    end else if(T1374) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1354) begin
      reqDone_6 <= 1'h0;
    end else if(T1352) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1332) begin
      reqDone_6 <= 1'h0;
    end else if(T1330) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1310) begin
      reqDone_6 <= 1'h0;
    end else if(T1308) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1288) begin
      reqDone_6 <= 1'h0;
    end else if(T1286) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1266) begin
      reqDone_6 <= 1'h0;
    end else if(T1264) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1244) begin
      reqDone_6 <= 1'h0;
    end else if(T1242) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1222) begin
      reqDone_6 <= 1'h0;
    end else if(T1220) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1200) begin
      reqDone_6 <= 1'h0;
    end else if(T1198) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1178) begin
      reqDone_6 <= 1'h0;
    end else if(T1176) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1156) begin
      reqDone_6 <= 1'h0;
    end else if(T1154) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1134) begin
      reqDone_6 <= 1'h0;
    end else if(T1132) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1112) begin
      reqDone_6 <= 1'h0;
    end else if(T1110) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1090) begin
      reqDone_6 <= 1'h0;
    end else if(T1088) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T1068) begin
      reqDone_6 <= 1'h0;
    end else if(T1066) begin
      reqDone_6 <= reqDoneWire_6;
    end else if(T86) begin
      reqDone_6 <= 1'h0;
    end
    if(reset) begin
      reqDone_5 <= 1'h0;
    end else if(T1484) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1464) begin
      reqDone_5 <= 1'h0;
    end else if(T1462) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1442) begin
      reqDone_5 <= 1'h0;
    end else if(T1440) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1420) begin
      reqDone_5 <= 1'h0;
    end else if(T1418) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1398) begin
      reqDone_5 <= 1'h0;
    end else if(T1396) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1376) begin
      reqDone_5 <= 1'h0;
    end else if(T1374) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1354) begin
      reqDone_5 <= 1'h0;
    end else if(T1352) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1332) begin
      reqDone_5 <= 1'h0;
    end else if(T1330) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1310) begin
      reqDone_5 <= 1'h0;
    end else if(T1308) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1288) begin
      reqDone_5 <= 1'h0;
    end else if(T1286) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1266) begin
      reqDone_5 <= 1'h0;
    end else if(T1264) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1244) begin
      reqDone_5 <= 1'h0;
    end else if(T1242) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1222) begin
      reqDone_5 <= 1'h0;
    end else if(T1220) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1200) begin
      reqDone_5 <= 1'h0;
    end else if(T1198) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1178) begin
      reqDone_5 <= 1'h0;
    end else if(T1176) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1156) begin
      reqDone_5 <= 1'h0;
    end else if(T1154) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1134) begin
      reqDone_5 <= 1'h0;
    end else if(T1132) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1112) begin
      reqDone_5 <= 1'h0;
    end else if(T1110) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1090) begin
      reqDone_5 <= 1'h0;
    end else if(T1088) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T1068) begin
      reqDone_5 <= 1'h0;
    end else if(T1066) begin
      reqDone_5 <= reqDoneWire_5;
    end else if(T86) begin
      reqDone_5 <= 1'h0;
    end
    if(reset) begin
      reqDone_4 <= 1'h0;
    end else if(T1484) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1464) begin
      reqDone_4 <= 1'h0;
    end else if(T1462) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1442) begin
      reqDone_4 <= 1'h0;
    end else if(T1440) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1420) begin
      reqDone_4 <= 1'h0;
    end else if(T1418) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1398) begin
      reqDone_4 <= 1'h0;
    end else if(T1396) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1376) begin
      reqDone_4 <= 1'h0;
    end else if(T1374) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1354) begin
      reqDone_4 <= 1'h0;
    end else if(T1352) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1332) begin
      reqDone_4 <= 1'h0;
    end else if(T1330) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1310) begin
      reqDone_4 <= 1'h0;
    end else if(T1308) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1288) begin
      reqDone_4 <= 1'h0;
    end else if(T1286) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1266) begin
      reqDone_4 <= 1'h0;
    end else if(T1264) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1244) begin
      reqDone_4 <= 1'h0;
    end else if(T1242) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1222) begin
      reqDone_4 <= 1'h0;
    end else if(T1220) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1200) begin
      reqDone_4 <= 1'h0;
    end else if(T1198) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1178) begin
      reqDone_4 <= 1'h0;
    end else if(T1176) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1156) begin
      reqDone_4 <= 1'h0;
    end else if(T1154) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1134) begin
      reqDone_4 <= 1'h0;
    end else if(T1132) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1112) begin
      reqDone_4 <= 1'h0;
    end else if(T1110) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1090) begin
      reqDone_4 <= 1'h0;
    end else if(T1088) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T1068) begin
      reqDone_4 <= 1'h0;
    end else if(T1066) begin
      reqDone_4 <= reqDoneWire_4;
    end else if(T86) begin
      reqDone_4 <= 1'h0;
    end
    if(reset) begin
      reqDone_3 <= 1'h0;
    end else if(T1484) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1464) begin
      reqDone_3 <= 1'h0;
    end else if(T1462) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1442) begin
      reqDone_3 <= 1'h0;
    end else if(T1440) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1420) begin
      reqDone_3 <= 1'h0;
    end else if(T1418) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1398) begin
      reqDone_3 <= 1'h0;
    end else if(T1396) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1376) begin
      reqDone_3 <= 1'h0;
    end else if(T1374) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1354) begin
      reqDone_3 <= 1'h0;
    end else if(T1352) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1332) begin
      reqDone_3 <= 1'h0;
    end else if(T1330) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1310) begin
      reqDone_3 <= 1'h0;
    end else if(T1308) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1288) begin
      reqDone_3 <= 1'h0;
    end else if(T1286) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1266) begin
      reqDone_3 <= 1'h0;
    end else if(T1264) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1244) begin
      reqDone_3 <= 1'h0;
    end else if(T1242) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1222) begin
      reqDone_3 <= 1'h0;
    end else if(T1220) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1200) begin
      reqDone_3 <= 1'h0;
    end else if(T1198) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1178) begin
      reqDone_3 <= 1'h0;
    end else if(T1176) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1156) begin
      reqDone_3 <= 1'h0;
    end else if(T1154) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1134) begin
      reqDone_3 <= 1'h0;
    end else if(T1132) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1112) begin
      reqDone_3 <= 1'h0;
    end else if(T1110) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1090) begin
      reqDone_3 <= 1'h0;
    end else if(T1088) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T1068) begin
      reqDone_3 <= 1'h0;
    end else if(T1066) begin
      reqDone_3 <= reqDoneWire_3;
    end else if(T86) begin
      reqDone_3 <= 1'h0;
    end
    if(reset) begin
      reqDone_2 <= 1'h0;
    end else if(T1484) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1464) begin
      reqDone_2 <= 1'h0;
    end else if(T1462) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1442) begin
      reqDone_2 <= 1'h0;
    end else if(T1440) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1420) begin
      reqDone_2 <= 1'h0;
    end else if(T1418) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1398) begin
      reqDone_2 <= 1'h0;
    end else if(T1396) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1376) begin
      reqDone_2 <= 1'h0;
    end else if(T1374) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1354) begin
      reqDone_2 <= 1'h0;
    end else if(T1352) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1332) begin
      reqDone_2 <= 1'h0;
    end else if(T1330) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1310) begin
      reqDone_2 <= 1'h0;
    end else if(T1308) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1288) begin
      reqDone_2 <= 1'h0;
    end else if(T1286) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1266) begin
      reqDone_2 <= 1'h0;
    end else if(T1264) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1244) begin
      reqDone_2 <= 1'h0;
    end else if(T1242) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1222) begin
      reqDone_2 <= 1'h0;
    end else if(T1220) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1200) begin
      reqDone_2 <= 1'h0;
    end else if(T1198) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1178) begin
      reqDone_2 <= 1'h0;
    end else if(T1176) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1156) begin
      reqDone_2 <= 1'h0;
    end else if(T1154) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1134) begin
      reqDone_2 <= 1'h0;
    end else if(T1132) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1112) begin
      reqDone_2 <= 1'h0;
    end else if(T1110) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1090) begin
      reqDone_2 <= 1'h0;
    end else if(T1088) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T1068) begin
      reqDone_2 <= 1'h0;
    end else if(T1066) begin
      reqDone_2 <= reqDoneWire_2;
    end else if(T86) begin
      reqDone_2 <= 1'h0;
    end
    if(reset) begin
      reqDone_1 <= 1'h0;
    end else if(T1484) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1464) begin
      reqDone_1 <= 1'h0;
    end else if(T1462) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1442) begin
      reqDone_1 <= 1'h0;
    end else if(T1440) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1420) begin
      reqDone_1 <= 1'h0;
    end else if(T1418) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1398) begin
      reqDone_1 <= 1'h0;
    end else if(T1396) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1376) begin
      reqDone_1 <= 1'h0;
    end else if(T1374) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1354) begin
      reqDone_1 <= 1'h0;
    end else if(T1352) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1332) begin
      reqDone_1 <= 1'h0;
    end else if(T1330) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1310) begin
      reqDone_1 <= 1'h0;
    end else if(T1308) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1288) begin
      reqDone_1 <= 1'h0;
    end else if(T1286) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1266) begin
      reqDone_1 <= 1'h0;
    end else if(T1264) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1244) begin
      reqDone_1 <= 1'h0;
    end else if(T1242) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1222) begin
      reqDone_1 <= 1'h0;
    end else if(T1220) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1200) begin
      reqDone_1 <= 1'h0;
    end else if(T1198) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1178) begin
      reqDone_1 <= 1'h0;
    end else if(T1176) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1156) begin
      reqDone_1 <= 1'h0;
    end else if(T1154) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1134) begin
      reqDone_1 <= 1'h0;
    end else if(T1132) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1112) begin
      reqDone_1 <= 1'h0;
    end else if(T1110) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1090) begin
      reqDone_1 <= 1'h0;
    end else if(T1088) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T1068) begin
      reqDone_1 <= 1'h0;
    end else if(T1066) begin
      reqDone_1 <= reqDoneWire_1;
    end else if(T86) begin
      reqDone_1 <= 1'h0;
    end
    seqMemAddr <= T1676;
    epilogueSpill <= T1679;
    if(reset) begin
      iterCount <= 32'h0;
    end else if(T1599) begin
      iterCount <= T1683;
    end
    if(reset) begin
      currentIter <= 32'h0;
    end else if(T1590) begin
      currentIter <= T1606;
    end else if(T1549) begin
      currentIter <= 32'h0;
    end
  end
endmodule

module customReg_4(input clk,
    input [57:0] io_inData,
    output[57:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [8:0] io_readAddr,
    input [8:0] io_writeAddr
);

  wire[57:0] T0;
  reg [57:0] ram [511:0];
  wire[57:0] T1;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 512; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];

  always @(posedge clk) begin
    if (io_writeEn)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module memConfig_10(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[8:0] io_memAddr,
    output[57:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[57:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[8:0] T87;
  reg [8:0] memAddr;
  wire[8:0] T97;
  wire[8:0] T88;
  wire[8:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h12;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h12;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h12;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h12;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[6'h39:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 9'h0;
  assign T97 = reset ? 9'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 9'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 9'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module fabOutSeqDP(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input [8:0] io_seqMemAddr,
    input  io_seqMemAddrValid,
    input [31:0] io_fabOut,
    input  io_fabOutValid,
    output io_fabOutRdy,
    output[31:0] io_fabOutStore,
    output io_fabOutStoreValid,
    input  io_fabOutStoreRdy,
    output[87:0] io_fabOutLoc,
    output io_fabOutLocValid,
    input  io_fabOutLocRdy,
    output io_seqProceed,
    output io_rst,
    output io_outLocValid
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  outDestLocal;
  wire T53;
  wire T5;
  wire T6;
  reg  outDestStore;
  wire T54;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire[57:0] nextSeq;
  wire[57:0] T14;
  wire T15;
  wire getNextSeq;
  wire T16;
  wire T17;
  reg  fabOutLocStrgValid;
  wire T55;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire seqDone;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg [87:0] fabOutLocStrg;
  wire[87:0] T56;
  wire[87:0] T48;
  wire[87:0] T49;
  wire[31:0] localStoreData;
  wire[55:0] bankInfo;
  wire[55:0] T50;
  wire[55:0] T51;
  wire[55:0] T52;
  wire[57:0] fabOutSeqMem_io_outData;
  wire fabOutSeqMemConfig_io_rst;
  wire[31:0] outStoreFifo_io_deqData;
  wire outStoreFifo_io_enqRdy;
  wire outStoreFifo_io_deqValid;
  wire[31:0] outLocalFifo_io_deqData;
  wire outLocalFifo_io_enqRdy;
  wire outLocalFifo_io_deqValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDestLocal = {1{$random}};
    outDestStore = {1{$random}};
    fabOutLocStrgValid = {1{$random}};
    fabOutLocStrg = {3{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = fabOutSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1 = T8 ? 1'h0 : T2;
  assign T2 = T3 ? io_fabOutValid : 1'h0;
  assign T3 = T6 & T4;
  assign T4 = outDestLocal & outLocalFifo_io_enqRdy;
  assign T53 = reset ? 1'h0 : T5;
  assign T5 = fabOutSeqMemConfig_io_rst ? 1'h0 : outDestLocal;
  assign T6 = outDestLocal | outDestStore;
  assign T54 = reset ? 1'h0 : T7;
  assign T7 = fabOutSeqMemConfig_io_rst ? 1'h0 : outDestStore;
  assign T8 = T6 & T9;
  assign T9 = T4 ^ 1'h1;
  assign T10 = T23 ? 1'h0 : T11;
  assign T11 = T12 ? 1'h1 : 1'h0;
  assign T12 = outLocalFifo_io_deqValid & T13;
  assign T13 = nextSeq[6'h38:6'h38];
  assign nextSeq = T14;
  assign T14 = T15 ? fabOutSeqMem_io_outData : 58'h0;
  assign T15 = T22 | getNextSeq;
  assign getNextSeq = T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = fabOutLocStrgValid & io_fabOutLocRdy;
  assign T55 = reset ? 1'h0 : T18;
  assign T18 = T17 ? 1'h0 : T19;
  assign T19 = outLocalFifo_io_deqValid ? 1'h1 : T20;
  assign T20 = fabOutSeqMemConfig_io_rst ? 1'h0 : fabOutLocStrgValid;
  assign T21 = T17 ^ 1'h1;
  assign T22 = ~ fabOutLocStrgValid;
  assign T23 = outLocalFifo_io_deqValid & T24;
  assign T24 = T13 ^ 1'h1;
  assign T25 = fabOutSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T26 = T30 ? 1'h0 : T27;
  assign T27 = T28 ? io_fabOutValid : 1'h0;
  assign T28 = T6 & T29;
  assign T29 = outDestStore & outStoreFifo_io_enqRdy;
  assign T30 = T6 & T31;
  assign T31 = T29 ^ 1'h1;
  assign io_outLocValid = outDestLocal;
  assign io_rst = fabOutSeqMemConfig_io_rst;
  assign io_seqProceed = T32;
  assign T32 = seqDone ? 1'h1 : 1'h0;
  assign seqDone = T33;
  assign T33 = T46 ? 1'h0 : T34;
  assign T34 = outLocalFifo_io_deqValid ? 1'h1 : T35;
  assign T35 = T43 ? 1'h1 : T36;
  assign T36 = T39 ? 1'h0 : T37;
  assign T37 = T15 & T38;
  assign T38 = ~ outDestLocal;
  assign T39 = T15 & T40;
  assign T40 = T42 & T41;
  assign T41 = nextSeq[6'h39:6'h39];
  assign T42 = T38 ^ 1'h1;
  assign T43 = T15 & T44;
  assign T44 = T45 ^ 1'h1;
  assign T45 = T38 | T41;
  assign T46 = outLocalFifo_io_deqValid ^ 1'h1;
  assign io_fabOutLocValid = T47;
  assign T47 = T17 ? fabOutLocStrgValid : 1'h0;
  assign io_fabOutLoc = fabOutLocStrg;
  assign T56 = reset ? 88'h0 : T48;
  assign T48 = outLocalFifo_io_deqValid ? T49 : fabOutLocStrg;
  assign T49 = {bankInfo, localStoreData};
  assign localStoreData = outLocalFifo_io_deqData;
  assign bankInfo = T50;
  assign T50 = T46 ? 56'h0 : T51;
  assign T51 = outLocalFifo_io_deqValid ? T52 : 56'h0;
  assign T52 = nextSeq[6'h37:1'h0];
  assign io_fabOutStoreValid = outStoreFifo_io_deqValid;
  assign io_fabOutStore = outStoreFifo_io_deqData;
  customReg_4 fabOutSeqMem(.clk(clk),
       //.io_inData(  )
       .io_outData( fabOutSeqMem_io_outData ),
       .io_readEn( io_seqMemAddrValid ),
       //.io_writeEn(  )
       .io_readAddr( io_seqMemAddr )
       //.io_writeAddr(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqMem.io_inData = {2{$random}};
    assign fabOutSeqMem.io_writeEn = {1{$random}};
    assign fabOutSeqMem.io_writeAddr = {1{$random}};
// synthesis translate_on
`endif
  memConfig_10 fabOutSeqMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       //.io_memAddr(  )
       //.io_memData(  )
       //.io_memOutValid(  )
       .io_rst( fabOutSeqMemConfig_io_rst )
  );
  fifo_1 outStoreFifo(.clk(clk), .reset(reset),
       .io_enqData( io_fabOut ),
       .io_deqData( outStoreFifo_io_deqData ),
       .io_enqRdy( outStoreFifo_io_enqRdy ),
       .io_deqRdy( io_fabOutStoreRdy ),
       .io_enqValid( T26 ),
       .io_deqValid( outStoreFifo_io_deqValid ),
       .io_rst( T25 )
  );
  fifo_1 outLocalFifo(.clk(clk), .reset(reset),
       .io_enqData( io_fabOut ),
       .io_deqData( outLocalFifo_io_deqData ),
       .io_enqRdy( outLocalFifo_io_enqRdy ),
       .io_deqRdy( T10 ),
       .io_enqValid( T1 ),
       .io_deqValid( outLocalFifo_io_deqValid ),
       .io_rst( T0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      outDestLocal <= 1'h0;
    end else if(fabOutSeqMemConfig_io_rst) begin
      outDestLocal <= 1'h0;
    end
    if(reset) begin
      outDestStore <= 1'h0;
    end else if(fabOutSeqMemConfig_io_rst) begin
      outDestStore <= 1'h0;
    end
    if(reset) begin
      fabOutLocStrgValid <= 1'h0;
    end else if(T17) begin
      fabOutLocStrgValid <= 1'h0;
    end else if(outLocalFifo_io_deqValid) begin
      fabOutLocStrgValid <= 1'h1;
    end else if(fabOutSeqMemConfig_io_rst) begin
      fabOutLocStrgValid <= 1'h0;
    end
    if(reset) begin
      fabOutLocStrg <= 88'h0;
    end else if(outLocalFifo_io_deqValid) begin
      fabOutLocStrg <= T49;
    end
  end
endmodule

module fabOutSeq(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input [31:0] io_fabOut_19,
    input [31:0] io_fabOut_18,
    input [31:0] io_fabOut_17,
    input [31:0] io_fabOut_16,
    input [31:0] io_fabOut_15,
    input [31:0] io_fabOut_14,
    input [31:0] io_fabOut_13,
    input [31:0] io_fabOut_12,
    input [31:0] io_fabOut_11,
    input [31:0] io_fabOut_10,
    input [31:0] io_fabOut_9,
    input [31:0] io_fabOut_8,
    input [31:0] io_fabOut_7,
    input [31:0] io_fabOut_6,
    input [31:0] io_fabOut_5,
    input [31:0] io_fabOut_4,
    input [31:0] io_fabOut_3,
    input [31:0] io_fabOut_2,
    input [31:0] io_fabOut_1,
    input [31:0] io_fabOut_0,
    input  io_fabOutValid_19,
    input  io_fabOutValid_18,
    input  io_fabOutValid_17,
    input  io_fabOutValid_16,
    input  io_fabOutValid_15,
    input  io_fabOutValid_14,
    input  io_fabOutValid_13,
    input  io_fabOutValid_12,
    input  io_fabOutValid_11,
    input  io_fabOutValid_10,
    input  io_fabOutValid_9,
    input  io_fabOutValid_8,
    input  io_fabOutValid_7,
    input  io_fabOutValid_6,
    input  io_fabOutValid_5,
    input  io_fabOutValid_4,
    input  io_fabOutValid_3,
    input  io_fabOutValid_2,
    input  io_fabOutValid_1,
    input  io_fabOutValid_0,
    output io_fabOutRdy_19,
    output io_fabOutRdy_18,
    output io_fabOutRdy_17,
    output io_fabOutRdy_16,
    output io_fabOutRdy_15,
    output io_fabOutRdy_14,
    output io_fabOutRdy_13,
    output io_fabOutRdy_12,
    output io_fabOutRdy_11,
    output io_fabOutRdy_10,
    output io_fabOutRdy_9,
    output io_fabOutRdy_8,
    output io_fabOutRdy_7,
    output io_fabOutRdy_6,
    output io_fabOutRdy_5,
    output io_fabOutRdy_4,
    output io_fabOutRdy_3,
    output io_fabOutRdy_2,
    output io_fabOutRdy_1,
    output io_fabOutRdy_0,
    output[31:0] io_fabOutStore_19,
    output[31:0] io_fabOutStore_18,
    output[31:0] io_fabOutStore_17,
    output[31:0] io_fabOutStore_16,
    output[31:0] io_fabOutStore_15,
    output[31:0] io_fabOutStore_14,
    output[31:0] io_fabOutStore_13,
    output[31:0] io_fabOutStore_12,
    output[31:0] io_fabOutStore_11,
    output[31:0] io_fabOutStore_10,
    output[31:0] io_fabOutStore_9,
    output[31:0] io_fabOutStore_8,
    output[31:0] io_fabOutStore_7,
    output[31:0] io_fabOutStore_6,
    output[31:0] io_fabOutStore_5,
    output[31:0] io_fabOutStore_4,
    output[31:0] io_fabOutStore_3,
    output[31:0] io_fabOutStore_2,
    output[31:0] io_fabOutStore_1,
    output[31:0] io_fabOutStore_0,
    output io_fabOutStoreValid_19,
    output io_fabOutStoreValid_18,
    output io_fabOutStoreValid_17,
    output io_fabOutStoreValid_16,
    output io_fabOutStoreValid_15,
    output io_fabOutStoreValid_14,
    output io_fabOutStoreValid_13,
    output io_fabOutStoreValid_12,
    output io_fabOutStoreValid_11,
    output io_fabOutStoreValid_10,
    output io_fabOutStoreValid_9,
    output io_fabOutStoreValid_8,
    output io_fabOutStoreValid_7,
    output io_fabOutStoreValid_6,
    output io_fabOutStoreValid_5,
    output io_fabOutStoreValid_4,
    output io_fabOutStoreValid_3,
    output io_fabOutStoreValid_2,
    output io_fabOutStoreValid_1,
    output io_fabOutStoreValid_0,
    input  io_fabOutStoreRdy_19,
    input  io_fabOutStoreRdy_18,
    input  io_fabOutStoreRdy_17,
    input  io_fabOutStoreRdy_16,
    input  io_fabOutStoreRdy_15,
    input  io_fabOutStoreRdy_14,
    input  io_fabOutStoreRdy_13,
    input  io_fabOutStoreRdy_12,
    input  io_fabOutStoreRdy_11,
    input  io_fabOutStoreRdy_10,
    input  io_fabOutStoreRdy_9,
    input  io_fabOutStoreRdy_8,
    input  io_fabOutStoreRdy_7,
    input  io_fabOutStoreRdy_6,
    input  io_fabOutStoreRdy_5,
    input  io_fabOutStoreRdy_4,
    input  io_fabOutStoreRdy_3,
    input  io_fabOutStoreRdy_2,
    input  io_fabOutStoreRdy_1,
    input  io_fabOutStoreRdy_0,
    output[87:0] io_fabOutLoc_19,
    output[87:0] io_fabOutLoc_18,
    output[87:0] io_fabOutLoc_17,
    output[87:0] io_fabOutLoc_16,
    output[87:0] io_fabOutLoc_15,
    output[87:0] io_fabOutLoc_14,
    output[87:0] io_fabOutLoc_13,
    output[87:0] io_fabOutLoc_12,
    output[87:0] io_fabOutLoc_11,
    output[87:0] io_fabOutLoc_10,
    output[87:0] io_fabOutLoc_9,
    output[87:0] io_fabOutLoc_8,
    output[87:0] io_fabOutLoc_7,
    output[87:0] io_fabOutLoc_6,
    output[87:0] io_fabOutLoc_5,
    output[87:0] io_fabOutLoc_4,
    output[87:0] io_fabOutLoc_3,
    output[87:0] io_fabOutLoc_2,
    output[87:0] io_fabOutLoc_1,
    output[87:0] io_fabOutLoc_0,
    output io_fabOutLocValid_19,
    output io_fabOutLocValid_18,
    output io_fabOutLocValid_17,
    output io_fabOutLocValid_16,
    output io_fabOutLocValid_15,
    output io_fabOutLocValid_14,
    output io_fabOutLocValid_13,
    output io_fabOutLocValid_12,
    output io_fabOutLocValid_11,
    output io_fabOutLocValid_10,
    output io_fabOutLocValid_9,
    output io_fabOutLocValid_8,
    output io_fabOutLocValid_7,
    output io_fabOutLocValid_6,
    output io_fabOutLocValid_5,
    output io_fabOutLocValid_4,
    output io_fabOutLocValid_3,
    output io_fabOutLocValid_2,
    output io_fabOutLocValid_1,
    output io_fabOutLocValid_0,
    input  io_fabOutLocRdy_19,
    input  io_fabOutLocRdy_18,
    input  io_fabOutLocRdy_17,
    input  io_fabOutLocRdy_16,
    input  io_fabOutLocRdy_15,
    input  io_fabOutLocRdy_14,
    input  io_fabOutLocRdy_13,
    input  io_fabOutLocRdy_12,
    input  io_fabOutLocRdy_11,
    input  io_fabOutLocRdy_10,
    input  io_fabOutLocRdy_9,
    input  io_fabOutLocRdy_8,
    input  io_fabOutLocRdy_7,
    input  io_fabOutLocRdy_6,
    input  io_fabOutLocRdy_5,
    input  io_fabOutLocRdy_4,
    input  io_fabOutLocRdy_3,
    input  io_fabOutLocRdy_2,
    input  io_fabOutLocRdy_1,
    input  io_fabOutLocRdy_0,
    output io_rst
);

  wire[8:0] fabOutCtrl_io_seqMemAddr_19;
  wire[8:0] fabOutCtrl_io_seqMemAddr_18;
  wire[8:0] fabOutCtrl_io_seqMemAddr_17;
  wire[8:0] fabOutCtrl_io_seqMemAddr_16;
  wire[8:0] fabOutCtrl_io_seqMemAddr_15;
  wire[8:0] fabOutCtrl_io_seqMemAddr_14;
  wire[8:0] fabOutCtrl_io_seqMemAddr_13;
  wire[8:0] fabOutCtrl_io_seqMemAddr_12;
  wire[8:0] fabOutCtrl_io_seqMemAddr_11;
  wire[8:0] fabOutCtrl_io_seqMemAddr_10;
  wire[8:0] fabOutCtrl_io_seqMemAddr_9;
  wire[8:0] fabOutCtrl_io_seqMemAddr_8;
  wire[8:0] fabOutCtrl_io_seqMemAddr_7;
  wire[8:0] fabOutCtrl_io_seqMemAddr_6;
  wire[8:0] fabOutCtrl_io_seqMemAddr_5;
  wire[8:0] fabOutCtrl_io_seqMemAddr_4;
  wire[8:0] fabOutCtrl_io_seqMemAddr_3;
  wire[8:0] fabOutCtrl_io_seqMemAddr_2;
  wire[8:0] fabOutCtrl_io_seqMemAddr_1;
  wire[8:0] fabOutCtrl_io_seqMemAddr_0;
  wire fabOutCtrl_io_seqMemAddrValid_19;
  wire fabOutCtrl_io_seqMemAddrValid_18;
  wire fabOutCtrl_io_seqMemAddrValid_17;
  wire fabOutCtrl_io_seqMemAddrValid_16;
  wire fabOutCtrl_io_seqMemAddrValid_15;
  wire fabOutCtrl_io_seqMemAddrValid_14;
  wire fabOutCtrl_io_seqMemAddrValid_13;
  wire fabOutCtrl_io_seqMemAddrValid_12;
  wire fabOutCtrl_io_seqMemAddrValid_11;
  wire fabOutCtrl_io_seqMemAddrValid_10;
  wire fabOutCtrl_io_seqMemAddrValid_9;
  wire fabOutCtrl_io_seqMemAddrValid_8;
  wire fabOutCtrl_io_seqMemAddrValid_7;
  wire fabOutCtrl_io_seqMemAddrValid_6;
  wire fabOutCtrl_io_seqMemAddrValid_5;
  wire fabOutCtrl_io_seqMemAddrValid_4;
  wire fabOutCtrl_io_seqMemAddrValid_3;
  wire fabOutCtrl_io_seqMemAddrValid_2;
  wire fabOutCtrl_io_seqMemAddrValid_1;
  wire fabOutCtrl_io_seqMemAddrValid_0;
  wire fabOutSeqDP_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_io_fabOutStore;
  wire fabOutSeqDP_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_io_fabOutLoc;
  wire fabOutSeqDP_io_fabOutLocValid;
  wire fabOutSeqDP_io_seqProceed;
  wire fabOutSeqDP_io_rst;
  wire fabOutSeqDP_io_outLocValid;
  wire fabOutSeqDP_1_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_1_io_fabOutStore;
  wire fabOutSeqDP_1_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_1_io_fabOutLoc;
  wire fabOutSeqDP_1_io_fabOutLocValid;
  wire fabOutSeqDP_1_io_seqProceed;
  wire fabOutSeqDP_1_io_outLocValid;
  wire fabOutSeqDP_2_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_2_io_fabOutStore;
  wire fabOutSeqDP_2_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_2_io_fabOutLoc;
  wire fabOutSeqDP_2_io_fabOutLocValid;
  wire fabOutSeqDP_2_io_seqProceed;
  wire fabOutSeqDP_2_io_outLocValid;
  wire fabOutSeqDP_3_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_3_io_fabOutStore;
  wire fabOutSeqDP_3_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_3_io_fabOutLoc;
  wire fabOutSeqDP_3_io_fabOutLocValid;
  wire fabOutSeqDP_3_io_seqProceed;
  wire fabOutSeqDP_3_io_outLocValid;
  wire fabOutSeqDP_4_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_4_io_fabOutStore;
  wire fabOutSeqDP_4_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_4_io_fabOutLoc;
  wire fabOutSeqDP_4_io_fabOutLocValid;
  wire fabOutSeqDP_4_io_seqProceed;
  wire fabOutSeqDP_4_io_outLocValid;
  wire fabOutSeqDP_5_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_5_io_fabOutStore;
  wire fabOutSeqDP_5_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_5_io_fabOutLoc;
  wire fabOutSeqDP_5_io_fabOutLocValid;
  wire fabOutSeqDP_5_io_seqProceed;
  wire fabOutSeqDP_5_io_outLocValid;
  wire fabOutSeqDP_6_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_6_io_fabOutStore;
  wire fabOutSeqDP_6_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_6_io_fabOutLoc;
  wire fabOutSeqDP_6_io_fabOutLocValid;
  wire fabOutSeqDP_6_io_seqProceed;
  wire fabOutSeqDP_6_io_outLocValid;
  wire fabOutSeqDP_7_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_7_io_fabOutStore;
  wire fabOutSeqDP_7_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_7_io_fabOutLoc;
  wire fabOutSeqDP_7_io_fabOutLocValid;
  wire fabOutSeqDP_7_io_seqProceed;
  wire fabOutSeqDP_7_io_outLocValid;
  wire fabOutSeqDP_8_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_8_io_fabOutStore;
  wire fabOutSeqDP_8_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_8_io_fabOutLoc;
  wire fabOutSeqDP_8_io_fabOutLocValid;
  wire fabOutSeqDP_8_io_seqProceed;
  wire fabOutSeqDP_8_io_outLocValid;
  wire fabOutSeqDP_9_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_9_io_fabOutStore;
  wire fabOutSeqDP_9_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_9_io_fabOutLoc;
  wire fabOutSeqDP_9_io_fabOutLocValid;
  wire fabOutSeqDP_9_io_seqProceed;
  wire fabOutSeqDP_9_io_outLocValid;
  wire fabOutSeqDP_10_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_10_io_fabOutStore;
  wire fabOutSeqDP_10_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_10_io_fabOutLoc;
  wire fabOutSeqDP_10_io_fabOutLocValid;
  wire fabOutSeqDP_10_io_seqProceed;
  wire fabOutSeqDP_10_io_outLocValid;
  wire fabOutSeqDP_11_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_11_io_fabOutStore;
  wire fabOutSeqDP_11_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_11_io_fabOutLoc;
  wire fabOutSeqDP_11_io_fabOutLocValid;
  wire fabOutSeqDP_11_io_seqProceed;
  wire fabOutSeqDP_11_io_outLocValid;
  wire fabOutSeqDP_12_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_12_io_fabOutStore;
  wire fabOutSeqDP_12_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_12_io_fabOutLoc;
  wire fabOutSeqDP_12_io_fabOutLocValid;
  wire fabOutSeqDP_12_io_seqProceed;
  wire fabOutSeqDP_12_io_outLocValid;
  wire fabOutSeqDP_13_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_13_io_fabOutStore;
  wire fabOutSeqDP_13_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_13_io_fabOutLoc;
  wire fabOutSeqDP_13_io_fabOutLocValid;
  wire fabOutSeqDP_13_io_seqProceed;
  wire fabOutSeqDP_13_io_outLocValid;
  wire fabOutSeqDP_14_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_14_io_fabOutStore;
  wire fabOutSeqDP_14_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_14_io_fabOutLoc;
  wire fabOutSeqDP_14_io_fabOutLocValid;
  wire fabOutSeqDP_14_io_seqProceed;
  wire fabOutSeqDP_14_io_outLocValid;
  wire fabOutSeqDP_15_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_15_io_fabOutStore;
  wire fabOutSeqDP_15_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_15_io_fabOutLoc;
  wire fabOutSeqDP_15_io_fabOutLocValid;
  wire fabOutSeqDP_15_io_seqProceed;
  wire fabOutSeqDP_15_io_outLocValid;
  wire fabOutSeqDP_16_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_16_io_fabOutStore;
  wire fabOutSeqDP_16_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_16_io_fabOutLoc;
  wire fabOutSeqDP_16_io_fabOutLocValid;
  wire fabOutSeqDP_16_io_seqProceed;
  wire fabOutSeqDP_16_io_outLocValid;
  wire fabOutSeqDP_17_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_17_io_fabOutStore;
  wire fabOutSeqDP_17_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_17_io_fabOutLoc;
  wire fabOutSeqDP_17_io_fabOutLocValid;
  wire fabOutSeqDP_17_io_seqProceed;
  wire fabOutSeqDP_17_io_outLocValid;
  wire fabOutSeqDP_18_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_18_io_fabOutStore;
  wire fabOutSeqDP_18_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_18_io_fabOutLoc;
  wire fabOutSeqDP_18_io_fabOutLocValid;
  wire fabOutSeqDP_18_io_seqProceed;
  wire fabOutSeqDP_18_io_outLocValid;
  wire fabOutSeqDP_19_io_fabOutRdy;
  wire[31:0] fabOutSeqDP_19_io_fabOutStore;
  wire fabOutSeqDP_19_io_fabOutStoreValid;
  wire[87:0] fabOutSeqDP_19_io_fabOutLoc;
  wire fabOutSeqDP_19_io_fabOutLocValid;
  wire fabOutSeqDP_19_io_seqProceed;
  wire fabOutSeqDP_19_io_outLocValid;


  assign io_rst = fabOutSeqDP_io_rst;
  assign io_fabOutLocValid_0 = fabOutSeqDP_io_fabOutLocValid;
  assign io_fabOutLocValid_1 = fabOutSeqDP_1_io_fabOutLocValid;
  assign io_fabOutLocValid_2 = fabOutSeqDP_2_io_fabOutLocValid;
  assign io_fabOutLocValid_3 = fabOutSeqDP_3_io_fabOutLocValid;
  assign io_fabOutLocValid_4 = fabOutSeqDP_4_io_fabOutLocValid;
  assign io_fabOutLocValid_5 = fabOutSeqDP_5_io_fabOutLocValid;
  assign io_fabOutLocValid_6 = fabOutSeqDP_6_io_fabOutLocValid;
  assign io_fabOutLocValid_7 = fabOutSeqDP_7_io_fabOutLocValid;
  assign io_fabOutLocValid_8 = fabOutSeqDP_8_io_fabOutLocValid;
  assign io_fabOutLocValid_9 = fabOutSeqDP_9_io_fabOutLocValid;
  assign io_fabOutLocValid_10 = fabOutSeqDP_10_io_fabOutLocValid;
  assign io_fabOutLocValid_11 = fabOutSeqDP_11_io_fabOutLocValid;
  assign io_fabOutLocValid_12 = fabOutSeqDP_12_io_fabOutLocValid;
  assign io_fabOutLocValid_13 = fabOutSeqDP_13_io_fabOutLocValid;
  assign io_fabOutLocValid_14 = fabOutSeqDP_14_io_fabOutLocValid;
  assign io_fabOutLocValid_15 = fabOutSeqDP_15_io_fabOutLocValid;
  assign io_fabOutLocValid_16 = fabOutSeqDP_16_io_fabOutLocValid;
  assign io_fabOutLocValid_17 = fabOutSeqDP_17_io_fabOutLocValid;
  assign io_fabOutLocValid_18 = fabOutSeqDP_18_io_fabOutLocValid;
  assign io_fabOutLocValid_19 = fabOutSeqDP_19_io_fabOutLocValid;
  assign io_fabOutLoc_0 = fabOutSeqDP_io_fabOutLoc;
  assign io_fabOutLoc_1 = fabOutSeqDP_1_io_fabOutLoc;
  assign io_fabOutLoc_2 = fabOutSeqDP_2_io_fabOutLoc;
  assign io_fabOutLoc_3 = fabOutSeqDP_3_io_fabOutLoc;
  assign io_fabOutLoc_4 = fabOutSeqDP_4_io_fabOutLoc;
  assign io_fabOutLoc_5 = fabOutSeqDP_5_io_fabOutLoc;
  assign io_fabOutLoc_6 = fabOutSeqDP_6_io_fabOutLoc;
  assign io_fabOutLoc_7 = fabOutSeqDP_7_io_fabOutLoc;
  assign io_fabOutLoc_8 = fabOutSeqDP_8_io_fabOutLoc;
  assign io_fabOutLoc_9 = fabOutSeqDP_9_io_fabOutLoc;
  assign io_fabOutLoc_10 = fabOutSeqDP_10_io_fabOutLoc;
  assign io_fabOutLoc_11 = fabOutSeqDP_11_io_fabOutLoc;
  assign io_fabOutLoc_12 = fabOutSeqDP_12_io_fabOutLoc;
  assign io_fabOutLoc_13 = fabOutSeqDP_13_io_fabOutLoc;
  assign io_fabOutLoc_14 = fabOutSeqDP_14_io_fabOutLoc;
  assign io_fabOutLoc_15 = fabOutSeqDP_15_io_fabOutLoc;
  assign io_fabOutLoc_16 = fabOutSeqDP_16_io_fabOutLoc;
  assign io_fabOutLoc_17 = fabOutSeqDP_17_io_fabOutLoc;
  assign io_fabOutLoc_18 = fabOutSeqDP_18_io_fabOutLoc;
  assign io_fabOutLoc_19 = fabOutSeqDP_19_io_fabOutLoc;
  assign io_fabOutStoreValid_0 = fabOutSeqDP_io_fabOutStoreValid;
  assign io_fabOutStoreValid_1 = fabOutSeqDP_1_io_fabOutStoreValid;
  assign io_fabOutStoreValid_2 = fabOutSeqDP_2_io_fabOutStoreValid;
  assign io_fabOutStoreValid_3 = fabOutSeqDP_3_io_fabOutStoreValid;
  assign io_fabOutStoreValid_4 = fabOutSeqDP_4_io_fabOutStoreValid;
  assign io_fabOutStoreValid_5 = fabOutSeqDP_5_io_fabOutStoreValid;
  assign io_fabOutStoreValid_6 = fabOutSeqDP_6_io_fabOutStoreValid;
  assign io_fabOutStoreValid_7 = fabOutSeqDP_7_io_fabOutStoreValid;
  assign io_fabOutStoreValid_8 = fabOutSeqDP_8_io_fabOutStoreValid;
  assign io_fabOutStoreValid_9 = fabOutSeqDP_9_io_fabOutStoreValid;
  assign io_fabOutStoreValid_10 = fabOutSeqDP_10_io_fabOutStoreValid;
  assign io_fabOutStoreValid_11 = fabOutSeqDP_11_io_fabOutStoreValid;
  assign io_fabOutStoreValid_12 = fabOutSeqDP_12_io_fabOutStoreValid;
  assign io_fabOutStoreValid_13 = fabOutSeqDP_13_io_fabOutStoreValid;
  assign io_fabOutStoreValid_14 = fabOutSeqDP_14_io_fabOutStoreValid;
  assign io_fabOutStoreValid_15 = fabOutSeqDP_15_io_fabOutStoreValid;
  assign io_fabOutStoreValid_16 = fabOutSeqDP_16_io_fabOutStoreValid;
  assign io_fabOutStoreValid_17 = fabOutSeqDP_17_io_fabOutStoreValid;
  assign io_fabOutStoreValid_18 = fabOutSeqDP_18_io_fabOutStoreValid;
  assign io_fabOutStoreValid_19 = fabOutSeqDP_19_io_fabOutStoreValid;
  assign io_fabOutStore_0 = fabOutSeqDP_io_fabOutStore;
  assign io_fabOutStore_1 = fabOutSeqDP_1_io_fabOutStore;
  assign io_fabOutStore_2 = fabOutSeqDP_2_io_fabOutStore;
  assign io_fabOutStore_3 = fabOutSeqDP_3_io_fabOutStore;
  assign io_fabOutStore_4 = fabOutSeqDP_4_io_fabOutStore;
  assign io_fabOutStore_5 = fabOutSeqDP_5_io_fabOutStore;
  assign io_fabOutStore_6 = fabOutSeqDP_6_io_fabOutStore;
  assign io_fabOutStore_7 = fabOutSeqDP_7_io_fabOutStore;
  assign io_fabOutStore_8 = fabOutSeqDP_8_io_fabOutStore;
  assign io_fabOutStore_9 = fabOutSeqDP_9_io_fabOutStore;
  assign io_fabOutStore_10 = fabOutSeqDP_10_io_fabOutStore;
  assign io_fabOutStore_11 = fabOutSeqDP_11_io_fabOutStore;
  assign io_fabOutStore_12 = fabOutSeqDP_12_io_fabOutStore;
  assign io_fabOutStore_13 = fabOutSeqDP_13_io_fabOutStore;
  assign io_fabOutStore_14 = fabOutSeqDP_14_io_fabOutStore;
  assign io_fabOutStore_15 = fabOutSeqDP_15_io_fabOutStore;
  assign io_fabOutStore_16 = fabOutSeqDP_16_io_fabOutStore;
  assign io_fabOutStore_17 = fabOutSeqDP_17_io_fabOutStore;
  assign io_fabOutStore_18 = fabOutSeqDP_18_io_fabOutStore;
  assign io_fabOutStore_19 = fabOutSeqDP_19_io_fabOutStore;
  assign io_fabOutRdy_0 = fabOutSeqDP_io_fabOutRdy;
  assign io_fabOutRdy_1 = fabOutSeqDP_1_io_fabOutRdy;
  assign io_fabOutRdy_2 = fabOutSeqDP_2_io_fabOutRdy;
  assign io_fabOutRdy_3 = fabOutSeqDP_3_io_fabOutRdy;
  assign io_fabOutRdy_4 = fabOutSeqDP_4_io_fabOutRdy;
  assign io_fabOutRdy_5 = fabOutSeqDP_5_io_fabOutRdy;
  assign io_fabOutRdy_6 = fabOutSeqDP_6_io_fabOutRdy;
  assign io_fabOutRdy_7 = fabOutSeqDP_7_io_fabOutRdy;
  assign io_fabOutRdy_8 = fabOutSeqDP_8_io_fabOutRdy;
  assign io_fabOutRdy_9 = fabOutSeqDP_9_io_fabOutRdy;
  assign io_fabOutRdy_10 = fabOutSeqDP_10_io_fabOutRdy;
  assign io_fabOutRdy_11 = fabOutSeqDP_11_io_fabOutRdy;
  assign io_fabOutRdy_12 = fabOutSeqDP_12_io_fabOutRdy;
  assign io_fabOutRdy_13 = fabOutSeqDP_13_io_fabOutRdy;
  assign io_fabOutRdy_14 = fabOutSeqDP_14_io_fabOutRdy;
  assign io_fabOutRdy_15 = fabOutSeqDP_15_io_fabOutRdy;
  assign io_fabOutRdy_16 = fabOutSeqDP_16_io_fabOutRdy;
  assign io_fabOutRdy_17 = fabOutSeqDP_17_io_fabOutRdy;
  assign io_fabOutRdy_18 = fabOutSeqDP_18_io_fabOutRdy;
  assign io_fabOutRdy_19 = fabOutSeqDP_19_io_fabOutRdy;
  fabOutSeqCtrl fabOutCtrl(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_outLocValid_19( fabOutSeqDP_19_io_outLocValid ),
       .io_outLocValid_18( fabOutSeqDP_18_io_outLocValid ),
       .io_outLocValid_17( fabOutSeqDP_17_io_outLocValid ),
       .io_outLocValid_16( fabOutSeqDP_16_io_outLocValid ),
       .io_outLocValid_15( fabOutSeqDP_15_io_outLocValid ),
       .io_outLocValid_14( fabOutSeqDP_14_io_outLocValid ),
       .io_outLocValid_13( fabOutSeqDP_13_io_outLocValid ),
       .io_outLocValid_12( fabOutSeqDP_12_io_outLocValid ),
       .io_outLocValid_11( fabOutSeqDP_11_io_outLocValid ),
       .io_outLocValid_10( fabOutSeqDP_10_io_outLocValid ),
       .io_outLocValid_9( fabOutSeqDP_9_io_outLocValid ),
       .io_outLocValid_8( fabOutSeqDP_8_io_outLocValid ),
       .io_outLocValid_7( fabOutSeqDP_7_io_outLocValid ),
       .io_outLocValid_6( fabOutSeqDP_6_io_outLocValid ),
       .io_outLocValid_5( fabOutSeqDP_5_io_outLocValid ),
       .io_outLocValid_4( fabOutSeqDP_4_io_outLocValid ),
       .io_outLocValid_3( fabOutSeqDP_3_io_outLocValid ),
       .io_outLocValid_2( fabOutSeqDP_2_io_outLocValid ),
       .io_outLocValid_1( fabOutSeqDP_1_io_outLocValid ),
       .io_outLocValid_0( fabOutSeqDP_io_outLocValid ),
       .io_seqMemAddr_19( fabOutCtrl_io_seqMemAddr_19 ),
       .io_seqMemAddr_18( fabOutCtrl_io_seqMemAddr_18 ),
       .io_seqMemAddr_17( fabOutCtrl_io_seqMemAddr_17 ),
       .io_seqMemAddr_16( fabOutCtrl_io_seqMemAddr_16 ),
       .io_seqMemAddr_15( fabOutCtrl_io_seqMemAddr_15 ),
       .io_seqMemAddr_14( fabOutCtrl_io_seqMemAddr_14 ),
       .io_seqMemAddr_13( fabOutCtrl_io_seqMemAddr_13 ),
       .io_seqMemAddr_12( fabOutCtrl_io_seqMemAddr_12 ),
       .io_seqMemAddr_11( fabOutCtrl_io_seqMemAddr_11 ),
       .io_seqMemAddr_10( fabOutCtrl_io_seqMemAddr_10 ),
       .io_seqMemAddr_9( fabOutCtrl_io_seqMemAddr_9 ),
       .io_seqMemAddr_8( fabOutCtrl_io_seqMemAddr_8 ),
       .io_seqMemAddr_7( fabOutCtrl_io_seqMemAddr_7 ),
       .io_seqMemAddr_6( fabOutCtrl_io_seqMemAddr_6 ),
       .io_seqMemAddr_5( fabOutCtrl_io_seqMemAddr_5 ),
       .io_seqMemAddr_4( fabOutCtrl_io_seqMemAddr_4 ),
       .io_seqMemAddr_3( fabOutCtrl_io_seqMemAddr_3 ),
       .io_seqMemAddr_2( fabOutCtrl_io_seqMemAddr_2 ),
       .io_seqMemAddr_1( fabOutCtrl_io_seqMemAddr_1 ),
       .io_seqMemAddr_0( fabOutCtrl_io_seqMemAddr_0 ),
       .io_seqMemAddrValid_19( fabOutCtrl_io_seqMemAddrValid_19 ),
       .io_seqMemAddrValid_18( fabOutCtrl_io_seqMemAddrValid_18 ),
       .io_seqMemAddrValid_17( fabOutCtrl_io_seqMemAddrValid_17 ),
       .io_seqMemAddrValid_16( fabOutCtrl_io_seqMemAddrValid_16 ),
       .io_seqMemAddrValid_15( fabOutCtrl_io_seqMemAddrValid_15 ),
       .io_seqMemAddrValid_14( fabOutCtrl_io_seqMemAddrValid_14 ),
       .io_seqMemAddrValid_13( fabOutCtrl_io_seqMemAddrValid_13 ),
       .io_seqMemAddrValid_12( fabOutCtrl_io_seqMemAddrValid_12 ),
       .io_seqMemAddrValid_11( fabOutCtrl_io_seqMemAddrValid_11 ),
       .io_seqMemAddrValid_10( fabOutCtrl_io_seqMemAddrValid_10 ),
       .io_seqMemAddrValid_9( fabOutCtrl_io_seqMemAddrValid_9 ),
       .io_seqMemAddrValid_8( fabOutCtrl_io_seqMemAddrValid_8 ),
       .io_seqMemAddrValid_7( fabOutCtrl_io_seqMemAddrValid_7 ),
       .io_seqMemAddrValid_6( fabOutCtrl_io_seqMemAddrValid_6 ),
       .io_seqMemAddrValid_5( fabOutCtrl_io_seqMemAddrValid_5 ),
       .io_seqMemAddrValid_4( fabOutCtrl_io_seqMemAddrValid_4 ),
       .io_seqMemAddrValid_3( fabOutCtrl_io_seqMemAddrValid_3 ),
       .io_seqMemAddrValid_2( fabOutCtrl_io_seqMemAddrValid_2 ),
       .io_seqMemAddrValid_1( fabOutCtrl_io_seqMemAddrValid_1 ),
       .io_seqMemAddrValid_0( fabOutCtrl_io_seqMemAddrValid_0 ),
       .io_seqProceed_19( fabOutSeqDP_19_io_seqProceed ),
       .io_seqProceed_18( fabOutSeqDP_18_io_seqProceed ),
       .io_seqProceed_17( fabOutSeqDP_17_io_seqProceed ),
       .io_seqProceed_16( fabOutSeqDP_16_io_seqProceed ),
       .io_seqProceed_15( fabOutSeqDP_15_io_seqProceed ),
       .io_seqProceed_14( fabOutSeqDP_14_io_seqProceed ),
       .io_seqProceed_13( fabOutSeqDP_13_io_seqProceed ),
       .io_seqProceed_12( fabOutSeqDP_12_io_seqProceed ),
       .io_seqProceed_11( fabOutSeqDP_11_io_seqProceed ),
       .io_seqProceed_10( fabOutSeqDP_10_io_seqProceed ),
       .io_seqProceed_9( fabOutSeqDP_9_io_seqProceed ),
       .io_seqProceed_8( fabOutSeqDP_8_io_seqProceed ),
       .io_seqProceed_7( fabOutSeqDP_7_io_seqProceed ),
       .io_seqProceed_6( fabOutSeqDP_6_io_seqProceed ),
       .io_seqProceed_5( fabOutSeqDP_5_io_seqProceed ),
       .io_seqProceed_4( fabOutSeqDP_4_io_seqProceed ),
       .io_seqProceed_3( fabOutSeqDP_3_io_seqProceed ),
       .io_seqProceed_2( fabOutSeqDP_2_io_seqProceed ),
       .io_seqProceed_1( fabOutSeqDP_1_io_seqProceed ),
       .io_seqProceed_0( fabOutSeqDP_io_seqProceed )
  );
  fabOutSeqDP fabOutSeqDP(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_0 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_0 ),
       .io_fabOut( io_fabOut_0 ),
       .io_fabOutValid( io_fabOutValid_0 ),
       .io_fabOutRdy( fabOutSeqDP_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_0 ),
       .io_fabOutLoc( fabOutSeqDP_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_0 ),
       .io_seqProceed( fabOutSeqDP_io_seqProceed ),
       .io_rst( fabOutSeqDP_io_rst ),
       .io_outLocValid( fabOutSeqDP_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_1(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_1 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_1 ),
       .io_fabOut( io_fabOut_1 ),
       .io_fabOutValid( io_fabOutValid_1 ),
       .io_fabOutRdy( fabOutSeqDP_1_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_1_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_1_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_1 ),
       .io_fabOutLoc( fabOutSeqDP_1_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_1_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_1 ),
       .io_seqProceed( fabOutSeqDP_1_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_1_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_1.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_2(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_2 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_2 ),
       .io_fabOut( io_fabOut_2 ),
       .io_fabOutValid( io_fabOutValid_2 ),
       .io_fabOutRdy( fabOutSeqDP_2_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_2_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_2_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_2 ),
       .io_fabOutLoc( fabOutSeqDP_2_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_2_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_2 ),
       .io_seqProceed( fabOutSeqDP_2_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_2_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_2.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_3(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_3 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_3 ),
       .io_fabOut( io_fabOut_3 ),
       .io_fabOutValid( io_fabOutValid_3 ),
       .io_fabOutRdy( fabOutSeqDP_3_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_3_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_3_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_3 ),
       .io_fabOutLoc( fabOutSeqDP_3_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_3_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_3 ),
       .io_seqProceed( fabOutSeqDP_3_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_3_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_3.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_4(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_4 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_4 ),
       .io_fabOut( io_fabOut_4 ),
       .io_fabOutValid( io_fabOutValid_4 ),
       .io_fabOutRdy( fabOutSeqDP_4_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_4_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_4_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_4 ),
       .io_fabOutLoc( fabOutSeqDP_4_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_4_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_4 ),
       .io_seqProceed( fabOutSeqDP_4_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_4_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_4.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_5(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_5 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_5 ),
       .io_fabOut( io_fabOut_5 ),
       .io_fabOutValid( io_fabOutValid_5 ),
       .io_fabOutRdy( fabOutSeqDP_5_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_5_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_5_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_5 ),
       .io_fabOutLoc( fabOutSeqDP_5_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_5_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_5 ),
       .io_seqProceed( fabOutSeqDP_5_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_5_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_5.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_6(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_6 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_6 ),
       .io_fabOut( io_fabOut_6 ),
       .io_fabOutValid( io_fabOutValid_6 ),
       .io_fabOutRdy( fabOutSeqDP_6_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_6_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_6_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_6 ),
       .io_fabOutLoc( fabOutSeqDP_6_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_6_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_6 ),
       .io_seqProceed( fabOutSeqDP_6_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_6_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_6.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_7(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_7 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_7 ),
       .io_fabOut( io_fabOut_7 ),
       .io_fabOutValid( io_fabOutValid_7 ),
       .io_fabOutRdy( fabOutSeqDP_7_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_7_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_7_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_7 ),
       .io_fabOutLoc( fabOutSeqDP_7_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_7_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_7 ),
       .io_seqProceed( fabOutSeqDP_7_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_7_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_7.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_8(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_8 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_8 ),
       .io_fabOut( io_fabOut_8 ),
       .io_fabOutValid( io_fabOutValid_8 ),
       .io_fabOutRdy( fabOutSeqDP_8_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_8_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_8_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_8 ),
       .io_fabOutLoc( fabOutSeqDP_8_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_8_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_8 ),
       .io_seqProceed( fabOutSeqDP_8_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_8_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_8.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_9(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_9 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_9 ),
       .io_fabOut( io_fabOut_9 ),
       .io_fabOutValid( io_fabOutValid_9 ),
       .io_fabOutRdy( fabOutSeqDP_9_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_9_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_9_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_9 ),
       .io_fabOutLoc( fabOutSeqDP_9_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_9_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_9 ),
       .io_seqProceed( fabOutSeqDP_9_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_9_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_9.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_10(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_10 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_10 ),
       .io_fabOut( io_fabOut_10 ),
       .io_fabOutValid( io_fabOutValid_10 ),
       .io_fabOutRdy( fabOutSeqDP_10_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_10_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_10_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_10 ),
       .io_fabOutLoc( fabOutSeqDP_10_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_10_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_10 ),
       .io_seqProceed( fabOutSeqDP_10_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_10_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_10.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_11(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_11 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_11 ),
       .io_fabOut( io_fabOut_11 ),
       .io_fabOutValid( io_fabOutValid_11 ),
       .io_fabOutRdy( fabOutSeqDP_11_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_11_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_11_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_11 ),
       .io_fabOutLoc( fabOutSeqDP_11_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_11_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_11 ),
       .io_seqProceed( fabOutSeqDP_11_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_11_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_11.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_12(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_12 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_12 ),
       .io_fabOut( io_fabOut_12 ),
       .io_fabOutValid( io_fabOutValid_12 ),
       .io_fabOutRdy( fabOutSeqDP_12_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_12_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_12_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_12 ),
       .io_fabOutLoc( fabOutSeqDP_12_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_12_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_12 ),
       .io_seqProceed( fabOutSeqDP_12_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_12_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_12.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_13(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_13 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_13 ),
       .io_fabOut( io_fabOut_13 ),
       .io_fabOutValid( io_fabOutValid_13 ),
       .io_fabOutRdy( fabOutSeqDP_13_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_13_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_13_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_13 ),
       .io_fabOutLoc( fabOutSeqDP_13_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_13_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_13 ),
       .io_seqProceed( fabOutSeqDP_13_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_13_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_13.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_14(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_14 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_14 ),
       .io_fabOut( io_fabOut_14 ),
       .io_fabOutValid( io_fabOutValid_14 ),
       .io_fabOutRdy( fabOutSeqDP_14_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_14_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_14_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_14 ),
       .io_fabOutLoc( fabOutSeqDP_14_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_14_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_14 ),
       .io_seqProceed( fabOutSeqDP_14_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_14_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_14.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_15(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_15 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_15 ),
       .io_fabOut( io_fabOut_15 ),
       .io_fabOutValid( io_fabOutValid_15 ),
       .io_fabOutRdy( fabOutSeqDP_15_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_15_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_15_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_15 ),
       .io_fabOutLoc( fabOutSeqDP_15_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_15_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_15 ),
       .io_seqProceed( fabOutSeqDP_15_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_15_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_15.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_16(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_16 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_16 ),
       .io_fabOut( io_fabOut_16 ),
       .io_fabOutValid( io_fabOutValid_16 ),
       .io_fabOutRdy( fabOutSeqDP_16_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_16_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_16_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_16 ),
       .io_fabOutLoc( fabOutSeqDP_16_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_16_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_16 ),
       .io_seqProceed( fabOutSeqDP_16_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_16_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_16.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_17(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_17 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_17 ),
       .io_fabOut( io_fabOut_17 ),
       .io_fabOutValid( io_fabOutValid_17 ),
       .io_fabOutRdy( fabOutSeqDP_17_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_17_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_17_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_17 ),
       .io_fabOutLoc( fabOutSeqDP_17_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_17_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_17 ),
       .io_seqProceed( fabOutSeqDP_17_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_17_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_17.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_18(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_18 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_18 ),
       .io_fabOut( io_fabOut_18 ),
       .io_fabOutValid( io_fabOutValid_18 ),
       .io_fabOutRdy( fabOutSeqDP_18_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_18_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_18_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_18 ),
       .io_fabOutLoc( fabOutSeqDP_18_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_18_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_18 ),
       .io_seqProceed( fabOutSeqDP_18_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_18_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_18.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
  fabOutSeqDP fabOutSeqDP_19(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_seqMemAddr( fabOutCtrl_io_seqMemAddr_19 ),
       .io_seqMemAddrValid( fabOutCtrl_io_seqMemAddrValid_19 ),
       .io_fabOut( io_fabOut_19 ),
       .io_fabOutValid( io_fabOutValid_19 ),
       .io_fabOutRdy( fabOutSeqDP_19_io_fabOutRdy ),
       .io_fabOutStore( fabOutSeqDP_19_io_fabOutStore ),
       .io_fabOutStoreValid( fabOutSeqDP_19_io_fabOutStoreValid ),
       .io_fabOutStoreRdy( io_fabOutStoreRdy_19 ),
       .io_fabOutLoc( fabOutSeqDP_19_io_fabOutLoc ),
       .io_fabOutLocValid( fabOutSeqDP_19_io_fabOutLocValid ),
       .io_fabOutLocRdy( io_fabOutLocRdy_19 ),
       .io_seqProceed( fabOutSeqDP_19_io_seqProceed ),
       //.io_rst(  )
       .io_outLocValid( fabOutSeqDP_19_io_outLocValid )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqDP_19.io_fabOutRdy = {1{$random}};
// synthesis translate_on
`endif
endmodule

module RRArbiter(input clk, input reset,
    input  io_request_19,
    input  io_request_18,
    input  io_request_17,
    input  io_request_16,
    input  io_request_15,
    input  io_request_14,
    input  io_request_13,
    input  io_request_12,
    input  io_request_11,
    input  io_request_10,
    input  io_request_9,
    input  io_request_8,
    input  io_request_7,
    input  io_request_6,
    input  io_request_5,
    input  io_request_4,
    input  io_request_3,
    input  io_request_2,
    input  io_request_1,
    input  io_request_0,
    output io_grant_19,
    output io_grant_18,
    output io_grant_17,
    output io_grant_16,
    output io_grant_15,
    output io_grant_14,
    output io_grant_13,
    output io_grant_12,
    output io_grant_11,
    output io_grant_10,
    output io_grant_9,
    output io_grant_8,
    output io_grant_7,
    output io_grant_6,
    output io_grant_5,
    output io_grant_4,
    output io_grant_3,
    output io_grant_2,
    output io_grant_1,
    output io_grant_0
);

  wire grant_0;
  wire T0;
  wire grantMasked_0;
  wire T1;
  wire T2;
  wire maskHihgerReq_0;
  wire requestMasked_0;
  wire T3;
  reg  pointerReg_0;
  wire T259;
  wire T4;
  wire T5;
  wire anyReqMasked;
  wire T6;
  wire requestMasked_19;
  wire T7;
  reg  pointerReg_19;
  wire T260;
  wire T8;
  wire T9;
  wire maskHihgerReq_19;
  wire T10;
  wire requestMasked_18;
  wire T11;
  reg  pointerReg_18;
  wire T261;
  wire T12;
  wire T13;
  wire unMaskHigherReq_18;
  wire T14;
  wire requestVec_17;
  wire unMaskHigherReq_17;
  wire T15;
  wire requestVec_16;
  wire unMaskHigherReq_16;
  wire T16;
  wire requestVec_15;
  wire unMaskHigherReq_15;
  wire T17;
  wire requestVec_14;
  wire unMaskHigherReq_14;
  wire T18;
  wire requestVec_13;
  wire unMaskHigherReq_13;
  wire T19;
  wire requestVec_12;
  wire unMaskHigherReq_12;
  wire T20;
  wire requestVec_11;
  wire unMaskHigherReq_11;
  wire T21;
  wire requestVec_10;
  wire unMaskHigherReq_10;
  wire T22;
  wire requestVec_9;
  wire unMaskHigherReq_9;
  wire T23;
  wire requestVec_8;
  wire unMaskHigherReq_8;
  wire T24;
  wire requestVec_7;
  wire unMaskHigherReq_7;
  wire T25;
  wire requestVec_6;
  wire unMaskHigherReq_6;
  wire T26;
  wire requestVec_5;
  wire unMaskHigherReq_5;
  wire T27;
  wire requestVec_4;
  wire unMaskHigherReq_4;
  wire T28;
  wire requestVec_3;
  wire unMaskHigherReq_3;
  wire T29;
  wire requestVec_2;
  wire unMaskHigherReq_2;
  wire T30;
  wire requestVec_1;
  wire unMaskHigherReq_1;
  wire T31;
  wire requestVec_18;
  wire maskHihgerReq_18;
  wire T32;
  wire requestMasked_17;
  wire T33;
  reg  pointerReg_17;
  wire T262;
  wire T34;
  wire T35;
  wire maskHihgerReq_17;
  wire T36;
  wire requestMasked_16;
  wire T37;
  reg  pointerReg_16;
  wire T263;
  wire T38;
  wire T39;
  wire maskHihgerReq_16;
  wire T40;
  wire requestMasked_15;
  wire T41;
  reg  pointerReg_15;
  wire T264;
  wire T42;
  wire T43;
  wire maskHihgerReq_15;
  wire T44;
  wire requestMasked_14;
  wire T45;
  reg  pointerReg_14;
  wire T265;
  wire T46;
  wire T47;
  wire maskHihgerReq_14;
  wire T48;
  wire requestMasked_13;
  wire T49;
  reg  pointerReg_13;
  wire T266;
  wire T50;
  wire T51;
  wire maskHihgerReq_13;
  wire T52;
  wire requestMasked_12;
  wire T53;
  reg  pointerReg_12;
  wire T267;
  wire T54;
  wire T55;
  wire maskHihgerReq_12;
  wire T56;
  wire requestMasked_11;
  wire T57;
  reg  pointerReg_11;
  wire T268;
  wire T58;
  wire T59;
  wire maskHihgerReq_11;
  wire T60;
  wire requestMasked_10;
  wire T61;
  reg  pointerReg_10;
  wire T269;
  wire T62;
  wire T63;
  wire maskHihgerReq_10;
  wire T64;
  wire requestMasked_9;
  wire T65;
  reg  pointerReg_9;
  wire T270;
  wire T66;
  wire T67;
  wire maskHihgerReq_9;
  wire T68;
  wire requestMasked_8;
  wire T69;
  reg  pointerReg_8;
  wire T271;
  wire T70;
  wire T71;
  wire maskHihgerReq_8;
  wire T72;
  wire requestMasked_7;
  wire T73;
  reg  pointerReg_7;
  wire T272;
  wire T74;
  wire T75;
  wire maskHihgerReq_7;
  wire T76;
  wire requestMasked_6;
  wire T77;
  reg  pointerReg_6;
  wire T273;
  wire T78;
  wire T79;
  wire maskHihgerReq_6;
  wire T80;
  wire requestMasked_5;
  wire T81;
  reg  pointerReg_5;
  wire T274;
  wire T82;
  wire T83;
  wire maskHihgerReq_5;
  wire T84;
  wire requestMasked_4;
  wire T85;
  reg  pointerReg_4;
  wire T275;
  wire T86;
  wire T87;
  wire maskHihgerReq_4;
  wire T88;
  wire requestMasked_3;
  wire T89;
  reg  pointerReg_3;
  wire T276;
  wire T90;
  wire T91;
  wire maskHihgerReq_3;
  wire T92;
  wire requestMasked_2;
  wire T93;
  reg  pointerReg_2;
  wire T277;
  wire T94;
  wire T95;
  wire maskHihgerReq_2;
  wire T96;
  wire requestMasked_1;
  wire T97;
  reg  pointerReg_1;
  wire T278;
  wire T98;
  wire T99;
  wire maskHihgerReq_1;
  wire T100;
  wire unMaskHigherReq_19;
  wire T101;
  wire requestVec_19;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire unMaskHigherReq_0;
  wire T120;
  wire requestAny;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire requestVec_0;
  wire T141;
  wire grantUnMasked_0;
  wire T142;
  wire T143;
  wire noReqMasked;
  wire T144;
  wire grant_1;
  wire T145;
  wire grantMasked_1;
  wire T146;
  wire T147;
  wire T148;
  wire grantUnMasked_1;
  wire T149;
  wire T150;
  wire grant_2;
  wire T151;
  wire grantMasked_2;
  wire T152;
  wire T153;
  wire T154;
  wire grantUnMasked_2;
  wire T155;
  wire T156;
  wire grant_3;
  wire T157;
  wire grantMasked_3;
  wire T158;
  wire T159;
  wire T160;
  wire grantUnMasked_3;
  wire T161;
  wire T162;
  wire grant_4;
  wire T163;
  wire grantMasked_4;
  wire T164;
  wire T165;
  wire T166;
  wire grantUnMasked_4;
  wire T167;
  wire T168;
  wire grant_5;
  wire T169;
  wire grantMasked_5;
  wire T170;
  wire T171;
  wire T172;
  wire grantUnMasked_5;
  wire T173;
  wire T174;
  wire grant_6;
  wire T175;
  wire grantMasked_6;
  wire T176;
  wire T177;
  wire T178;
  wire grantUnMasked_6;
  wire T179;
  wire T180;
  wire grant_7;
  wire T181;
  wire grantMasked_7;
  wire T182;
  wire T183;
  wire T184;
  wire grantUnMasked_7;
  wire T185;
  wire T186;
  wire grant_8;
  wire T187;
  wire grantMasked_8;
  wire T188;
  wire T189;
  wire T190;
  wire grantUnMasked_8;
  wire T191;
  wire T192;
  wire grant_9;
  wire T193;
  wire grantMasked_9;
  wire T194;
  wire T195;
  wire T196;
  wire grantUnMasked_9;
  wire T197;
  wire T198;
  wire grant_10;
  wire T199;
  wire grantMasked_10;
  wire T200;
  wire T201;
  wire T202;
  wire grantUnMasked_10;
  wire T203;
  wire T204;
  wire grant_11;
  wire T205;
  wire grantMasked_11;
  wire T206;
  wire T207;
  wire T208;
  wire grantUnMasked_11;
  wire T209;
  wire T210;
  wire grant_12;
  wire T211;
  wire grantMasked_12;
  wire T212;
  wire T213;
  wire T214;
  wire grantUnMasked_12;
  wire T215;
  wire T216;
  wire grant_13;
  wire T217;
  wire grantMasked_13;
  wire T218;
  wire T219;
  wire T220;
  wire grantUnMasked_13;
  wire T221;
  wire T222;
  wire grant_14;
  wire T223;
  wire grantMasked_14;
  wire T224;
  wire T225;
  wire T226;
  wire grantUnMasked_14;
  wire T227;
  wire T228;
  wire grant_15;
  wire T229;
  wire grantMasked_15;
  wire T230;
  wire T231;
  wire T232;
  wire grantUnMasked_15;
  wire T233;
  wire T234;
  wire grant_16;
  wire T235;
  wire grantMasked_16;
  wire T236;
  wire T237;
  wire T238;
  wire grantUnMasked_16;
  wire T239;
  wire T240;
  wire grant_17;
  wire T241;
  wire grantMasked_17;
  wire T242;
  wire T243;
  wire T244;
  wire grantUnMasked_17;
  wire T245;
  wire T246;
  wire grant_18;
  wire T247;
  wire grantMasked_18;
  wire T248;
  wire T249;
  wire T250;
  wire grantUnMasked_18;
  wire T251;
  wire T252;
  wire grant_19;
  wire T253;
  wire grantMasked_19;
  wire T254;
  wire T255;
  wire T256;
  wire grantUnMasked_19;
  wire T257;
  wire T258;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    pointerReg_0 = {1{$random}};
    pointerReg_19 = {1{$random}};
    pointerReg_18 = {1{$random}};
    pointerReg_17 = {1{$random}};
    pointerReg_16 = {1{$random}};
    pointerReg_15 = {1{$random}};
    pointerReg_14 = {1{$random}};
    pointerReg_13 = {1{$random}};
    pointerReg_12 = {1{$random}};
    pointerReg_11 = {1{$random}};
    pointerReg_10 = {1{$random}};
    pointerReg_9 = {1{$random}};
    pointerReg_8 = {1{$random}};
    pointerReg_7 = {1{$random}};
    pointerReg_6 = {1{$random}};
    pointerReg_5 = {1{$random}};
    pointerReg_4 = {1{$random}};
    pointerReg_3 = {1{$random}};
    pointerReg_2 = {1{$random}};
    pointerReg_1 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign maskHihgerReq_0 = {1{$random}};
  assign unMaskHigherReq_0 = {1{$random}};
// synthesis translate_on
`endif
  assign io_grant_0 = grant_0;
  assign grant_0 = T0;
  assign T0 = T141 | grantMasked_0;
  assign grantMasked_0 = T1;
  assign T1 = requestMasked_0 & T2;
  assign T2 = ~ maskHihgerReq_0;
  assign requestMasked_0 = T3;
  assign T3 = requestVec_0 & pointerReg_0;
  assign T259 = reset ? 1'h0 : T4;
  assign T4 = T120 ? unMaskHigherReq_0 : T5;
  assign T5 = anyReqMasked ? maskHihgerReq_0 : pointerReg_0;
  assign anyReqMasked = T6;
  assign T6 = T102 | requestMasked_19;
  assign requestMasked_19 = T7;
  assign T7 = requestVec_19 & pointerReg_19;
  assign T260 = reset ? 1'h0 : T8;
  assign T8 = T120 ? unMaskHigherReq_19 : T9;
  assign T9 = anyReqMasked ? maskHihgerReq_19 : pointerReg_19;
  assign maskHihgerReq_19 = T10;
  assign T10 = maskHihgerReq_18 | requestMasked_18;
  assign requestMasked_18 = T11;
  assign T11 = requestVec_18 & pointerReg_18;
  assign T261 = reset ? 1'h0 : T12;
  assign T12 = T120 ? unMaskHigherReq_18 : T13;
  assign T13 = anyReqMasked ? maskHihgerReq_18 : pointerReg_18;
  assign unMaskHigherReq_18 = T14;
  assign T14 = unMaskHigherReq_17 | requestVec_17;
  assign requestVec_17 = io_request_17;
  assign unMaskHigherReq_17 = T15;
  assign T15 = unMaskHigherReq_16 | requestVec_16;
  assign requestVec_16 = io_request_16;
  assign unMaskHigherReq_16 = T16;
  assign T16 = unMaskHigherReq_15 | requestVec_15;
  assign requestVec_15 = io_request_15;
  assign unMaskHigherReq_15 = T17;
  assign T17 = unMaskHigherReq_14 | requestVec_14;
  assign requestVec_14 = io_request_14;
  assign unMaskHigherReq_14 = T18;
  assign T18 = unMaskHigherReq_13 | requestVec_13;
  assign requestVec_13 = io_request_13;
  assign unMaskHigherReq_13 = T19;
  assign T19 = unMaskHigherReq_12 | requestVec_12;
  assign requestVec_12 = io_request_12;
  assign unMaskHigherReq_12 = T20;
  assign T20 = unMaskHigherReq_11 | requestVec_11;
  assign requestVec_11 = io_request_11;
  assign unMaskHigherReq_11 = T21;
  assign T21 = unMaskHigherReq_10 | requestVec_10;
  assign requestVec_10 = io_request_10;
  assign unMaskHigherReq_10 = T22;
  assign T22 = unMaskHigherReq_9 | requestVec_9;
  assign requestVec_9 = io_request_9;
  assign unMaskHigherReq_9 = T23;
  assign T23 = unMaskHigherReq_8 | requestVec_8;
  assign requestVec_8 = io_request_8;
  assign unMaskHigherReq_8 = T24;
  assign T24 = unMaskHigherReq_7 | requestVec_7;
  assign requestVec_7 = io_request_7;
  assign unMaskHigherReq_7 = T25;
  assign T25 = unMaskHigherReq_6 | requestVec_6;
  assign requestVec_6 = io_request_6;
  assign unMaskHigherReq_6 = T26;
  assign T26 = unMaskHigherReq_5 | requestVec_5;
  assign requestVec_5 = io_request_5;
  assign unMaskHigherReq_5 = T27;
  assign T27 = unMaskHigherReq_4 | requestVec_4;
  assign requestVec_4 = io_request_4;
  assign unMaskHigherReq_4 = T28;
  assign T28 = unMaskHigherReq_3 | requestVec_3;
  assign requestVec_3 = io_request_3;
  assign unMaskHigherReq_3 = T29;
  assign T29 = unMaskHigherReq_2 | requestVec_2;
  assign requestVec_2 = io_request_2;
  assign unMaskHigherReq_2 = T30;
  assign T30 = unMaskHigherReq_1 | requestVec_1;
  assign requestVec_1 = io_request_1;
  assign unMaskHigherReq_1 = T31;
  assign T31 = unMaskHigherReq_0 | requestVec_0;
  assign requestVec_18 = io_request_18;
  assign maskHihgerReq_18 = T32;
  assign T32 = maskHihgerReq_17 | requestMasked_17;
  assign requestMasked_17 = T33;
  assign T33 = requestVec_17 & pointerReg_17;
  assign T262 = reset ? 1'h0 : T34;
  assign T34 = T120 ? unMaskHigherReq_17 : T35;
  assign T35 = anyReqMasked ? maskHihgerReq_17 : pointerReg_17;
  assign maskHihgerReq_17 = T36;
  assign T36 = maskHihgerReq_16 | requestMasked_16;
  assign requestMasked_16 = T37;
  assign T37 = requestVec_16 & pointerReg_16;
  assign T263 = reset ? 1'h0 : T38;
  assign T38 = T120 ? unMaskHigherReq_16 : T39;
  assign T39 = anyReqMasked ? maskHihgerReq_16 : pointerReg_16;
  assign maskHihgerReq_16 = T40;
  assign T40 = maskHihgerReq_15 | requestMasked_15;
  assign requestMasked_15 = T41;
  assign T41 = requestVec_15 & pointerReg_15;
  assign T264 = reset ? 1'h0 : T42;
  assign T42 = T120 ? unMaskHigherReq_15 : T43;
  assign T43 = anyReqMasked ? maskHihgerReq_15 : pointerReg_15;
  assign maskHihgerReq_15 = T44;
  assign T44 = maskHihgerReq_14 | requestMasked_14;
  assign requestMasked_14 = T45;
  assign T45 = requestVec_14 & pointerReg_14;
  assign T265 = reset ? 1'h0 : T46;
  assign T46 = T120 ? unMaskHigherReq_14 : T47;
  assign T47 = anyReqMasked ? maskHihgerReq_14 : pointerReg_14;
  assign maskHihgerReq_14 = T48;
  assign T48 = maskHihgerReq_13 | requestMasked_13;
  assign requestMasked_13 = T49;
  assign T49 = requestVec_13 & pointerReg_13;
  assign T266 = reset ? 1'h0 : T50;
  assign T50 = T120 ? unMaskHigherReq_13 : T51;
  assign T51 = anyReqMasked ? maskHihgerReq_13 : pointerReg_13;
  assign maskHihgerReq_13 = T52;
  assign T52 = maskHihgerReq_12 | requestMasked_12;
  assign requestMasked_12 = T53;
  assign T53 = requestVec_12 & pointerReg_12;
  assign T267 = reset ? 1'h0 : T54;
  assign T54 = T120 ? unMaskHigherReq_12 : T55;
  assign T55 = anyReqMasked ? maskHihgerReq_12 : pointerReg_12;
  assign maskHihgerReq_12 = T56;
  assign T56 = maskHihgerReq_11 | requestMasked_11;
  assign requestMasked_11 = T57;
  assign T57 = requestVec_11 & pointerReg_11;
  assign T268 = reset ? 1'h0 : T58;
  assign T58 = T120 ? unMaskHigherReq_11 : T59;
  assign T59 = anyReqMasked ? maskHihgerReq_11 : pointerReg_11;
  assign maskHihgerReq_11 = T60;
  assign T60 = maskHihgerReq_10 | requestMasked_10;
  assign requestMasked_10 = T61;
  assign T61 = requestVec_10 & pointerReg_10;
  assign T269 = reset ? 1'h0 : T62;
  assign T62 = T120 ? unMaskHigherReq_10 : T63;
  assign T63 = anyReqMasked ? maskHihgerReq_10 : pointerReg_10;
  assign maskHihgerReq_10 = T64;
  assign T64 = maskHihgerReq_9 | requestMasked_9;
  assign requestMasked_9 = T65;
  assign T65 = requestVec_9 & pointerReg_9;
  assign T270 = reset ? 1'h0 : T66;
  assign T66 = T120 ? unMaskHigherReq_9 : T67;
  assign T67 = anyReqMasked ? maskHihgerReq_9 : pointerReg_9;
  assign maskHihgerReq_9 = T68;
  assign T68 = maskHihgerReq_8 | requestMasked_8;
  assign requestMasked_8 = T69;
  assign T69 = requestVec_8 & pointerReg_8;
  assign T271 = reset ? 1'h0 : T70;
  assign T70 = T120 ? unMaskHigherReq_8 : T71;
  assign T71 = anyReqMasked ? maskHihgerReq_8 : pointerReg_8;
  assign maskHihgerReq_8 = T72;
  assign T72 = maskHihgerReq_7 | requestMasked_7;
  assign requestMasked_7 = T73;
  assign T73 = requestVec_7 & pointerReg_7;
  assign T272 = reset ? 1'h0 : T74;
  assign T74 = T120 ? unMaskHigherReq_7 : T75;
  assign T75 = anyReqMasked ? maskHihgerReq_7 : pointerReg_7;
  assign maskHihgerReq_7 = T76;
  assign T76 = maskHihgerReq_6 | requestMasked_6;
  assign requestMasked_6 = T77;
  assign T77 = requestVec_6 & pointerReg_6;
  assign T273 = reset ? 1'h0 : T78;
  assign T78 = T120 ? unMaskHigherReq_6 : T79;
  assign T79 = anyReqMasked ? maskHihgerReq_6 : pointerReg_6;
  assign maskHihgerReq_6 = T80;
  assign T80 = maskHihgerReq_5 | requestMasked_5;
  assign requestMasked_5 = T81;
  assign T81 = requestVec_5 & pointerReg_5;
  assign T274 = reset ? 1'h0 : T82;
  assign T82 = T120 ? unMaskHigherReq_5 : T83;
  assign T83 = anyReqMasked ? maskHihgerReq_5 : pointerReg_5;
  assign maskHihgerReq_5 = T84;
  assign T84 = maskHihgerReq_4 | requestMasked_4;
  assign requestMasked_4 = T85;
  assign T85 = requestVec_4 & pointerReg_4;
  assign T275 = reset ? 1'h0 : T86;
  assign T86 = T120 ? unMaskHigherReq_4 : T87;
  assign T87 = anyReqMasked ? maskHihgerReq_4 : pointerReg_4;
  assign maskHihgerReq_4 = T88;
  assign T88 = maskHihgerReq_3 | requestMasked_3;
  assign requestMasked_3 = T89;
  assign T89 = requestVec_3 & pointerReg_3;
  assign T276 = reset ? 1'h0 : T90;
  assign T90 = T120 ? unMaskHigherReq_3 : T91;
  assign T91 = anyReqMasked ? maskHihgerReq_3 : pointerReg_3;
  assign maskHihgerReq_3 = T92;
  assign T92 = maskHihgerReq_2 | requestMasked_2;
  assign requestMasked_2 = T93;
  assign T93 = requestVec_2 & pointerReg_2;
  assign T277 = reset ? 1'h0 : T94;
  assign T94 = T120 ? unMaskHigherReq_2 : T95;
  assign T95 = anyReqMasked ? maskHihgerReq_2 : pointerReg_2;
  assign maskHihgerReq_2 = T96;
  assign T96 = maskHihgerReq_1 | requestMasked_1;
  assign requestMasked_1 = T97;
  assign T97 = requestVec_1 & pointerReg_1;
  assign T278 = reset ? 1'h0 : T98;
  assign T98 = T120 ? unMaskHigherReq_1 : T99;
  assign T99 = anyReqMasked ? maskHihgerReq_1 : pointerReg_1;
  assign maskHihgerReq_1 = T100;
  assign T100 = maskHihgerReq_0 | requestMasked_0;
  assign unMaskHigherReq_19 = T101;
  assign T101 = unMaskHigherReq_18 | requestVec_18;
  assign requestVec_19 = io_request_19;
  assign T102 = T103 | requestMasked_18;
  assign T103 = T104 | requestMasked_17;
  assign T104 = T105 | requestMasked_16;
  assign T105 = T106 | requestMasked_15;
  assign T106 = T107 | requestMasked_14;
  assign T107 = T108 | requestMasked_13;
  assign T108 = T109 | requestMasked_12;
  assign T109 = T110 | requestMasked_11;
  assign T110 = T111 | requestMasked_10;
  assign T111 = T112 | requestMasked_9;
  assign T112 = T113 | requestMasked_8;
  assign T113 = T114 | requestMasked_7;
  assign T114 = T115 | requestMasked_6;
  assign T115 = T116 | requestMasked_5;
  assign T116 = T117 | requestMasked_4;
  assign T117 = T118 | requestMasked_3;
  assign T118 = T119 | requestMasked_2;
  assign T119 = requestMasked_0 | requestMasked_1;
  assign T120 = T140 & requestAny;
  assign requestAny = T121;
  assign T121 = T122 | requestVec_19;
  assign T122 = T123 | requestVec_18;
  assign T123 = T124 | requestVec_17;
  assign T124 = T125 | requestVec_16;
  assign T125 = T126 | requestVec_15;
  assign T126 = T127 | requestVec_14;
  assign T127 = T128 | requestVec_13;
  assign T128 = T129 | requestVec_12;
  assign T129 = T130 | requestVec_11;
  assign T130 = T131 | requestVec_10;
  assign T131 = T132 | requestVec_9;
  assign T132 = T133 | requestVec_8;
  assign T133 = T134 | requestVec_7;
  assign T134 = T135 | requestVec_6;
  assign T135 = T136 | requestVec_5;
  assign T136 = T137 | requestVec_4;
  assign T137 = T138 | requestVec_3;
  assign T138 = T139 | requestVec_2;
  assign T139 = requestVec_0 | requestVec_1;
  assign T140 = anyReqMasked ^ 1'h1;
  assign requestVec_0 = io_request_0;
  assign T141 = noReqMasked & grantUnMasked_0;
  assign grantUnMasked_0 = T142;
  assign T142 = requestVec_0 & T143;
  assign T143 = ~ unMaskHigherReq_0;
  assign noReqMasked = T144;
  assign T144 = ~ anyReqMasked;
  assign io_grant_1 = grant_1;
  assign grant_1 = T145;
  assign T145 = T148 | grantMasked_1;
  assign grantMasked_1 = T146;
  assign T146 = requestMasked_1 & T147;
  assign T147 = ~ maskHihgerReq_1;
  assign T148 = noReqMasked & grantUnMasked_1;
  assign grantUnMasked_1 = T149;
  assign T149 = requestVec_1 & T150;
  assign T150 = ~ unMaskHigherReq_1;
  assign io_grant_2 = grant_2;
  assign grant_2 = T151;
  assign T151 = T154 | grantMasked_2;
  assign grantMasked_2 = T152;
  assign T152 = requestMasked_2 & T153;
  assign T153 = ~ maskHihgerReq_2;
  assign T154 = noReqMasked & grantUnMasked_2;
  assign grantUnMasked_2 = T155;
  assign T155 = requestVec_2 & T156;
  assign T156 = ~ unMaskHigherReq_2;
  assign io_grant_3 = grant_3;
  assign grant_3 = T157;
  assign T157 = T160 | grantMasked_3;
  assign grantMasked_3 = T158;
  assign T158 = requestMasked_3 & T159;
  assign T159 = ~ maskHihgerReq_3;
  assign T160 = noReqMasked & grantUnMasked_3;
  assign grantUnMasked_3 = T161;
  assign T161 = requestVec_3 & T162;
  assign T162 = ~ unMaskHigherReq_3;
  assign io_grant_4 = grant_4;
  assign grant_4 = T163;
  assign T163 = T166 | grantMasked_4;
  assign grantMasked_4 = T164;
  assign T164 = requestMasked_4 & T165;
  assign T165 = ~ maskHihgerReq_4;
  assign T166 = noReqMasked & grantUnMasked_4;
  assign grantUnMasked_4 = T167;
  assign T167 = requestVec_4 & T168;
  assign T168 = ~ unMaskHigherReq_4;
  assign io_grant_5 = grant_5;
  assign grant_5 = T169;
  assign T169 = T172 | grantMasked_5;
  assign grantMasked_5 = T170;
  assign T170 = requestMasked_5 & T171;
  assign T171 = ~ maskHihgerReq_5;
  assign T172 = noReqMasked & grantUnMasked_5;
  assign grantUnMasked_5 = T173;
  assign T173 = requestVec_5 & T174;
  assign T174 = ~ unMaskHigherReq_5;
  assign io_grant_6 = grant_6;
  assign grant_6 = T175;
  assign T175 = T178 | grantMasked_6;
  assign grantMasked_6 = T176;
  assign T176 = requestMasked_6 & T177;
  assign T177 = ~ maskHihgerReq_6;
  assign T178 = noReqMasked & grantUnMasked_6;
  assign grantUnMasked_6 = T179;
  assign T179 = requestVec_6 & T180;
  assign T180 = ~ unMaskHigherReq_6;
  assign io_grant_7 = grant_7;
  assign grant_7 = T181;
  assign T181 = T184 | grantMasked_7;
  assign grantMasked_7 = T182;
  assign T182 = requestMasked_7 & T183;
  assign T183 = ~ maskHihgerReq_7;
  assign T184 = noReqMasked & grantUnMasked_7;
  assign grantUnMasked_7 = T185;
  assign T185 = requestVec_7 & T186;
  assign T186 = ~ unMaskHigherReq_7;
  assign io_grant_8 = grant_8;
  assign grant_8 = T187;
  assign T187 = T190 | grantMasked_8;
  assign grantMasked_8 = T188;
  assign T188 = requestMasked_8 & T189;
  assign T189 = ~ maskHihgerReq_8;
  assign T190 = noReqMasked & grantUnMasked_8;
  assign grantUnMasked_8 = T191;
  assign T191 = requestVec_8 & T192;
  assign T192 = ~ unMaskHigherReq_8;
  assign io_grant_9 = grant_9;
  assign grant_9 = T193;
  assign T193 = T196 | grantMasked_9;
  assign grantMasked_9 = T194;
  assign T194 = requestMasked_9 & T195;
  assign T195 = ~ maskHihgerReq_9;
  assign T196 = noReqMasked & grantUnMasked_9;
  assign grantUnMasked_9 = T197;
  assign T197 = requestVec_9 & T198;
  assign T198 = ~ unMaskHigherReq_9;
  assign io_grant_10 = grant_10;
  assign grant_10 = T199;
  assign T199 = T202 | grantMasked_10;
  assign grantMasked_10 = T200;
  assign T200 = requestMasked_10 & T201;
  assign T201 = ~ maskHihgerReq_10;
  assign T202 = noReqMasked & grantUnMasked_10;
  assign grantUnMasked_10 = T203;
  assign T203 = requestVec_10 & T204;
  assign T204 = ~ unMaskHigherReq_10;
  assign io_grant_11 = grant_11;
  assign grant_11 = T205;
  assign T205 = T208 | grantMasked_11;
  assign grantMasked_11 = T206;
  assign T206 = requestMasked_11 & T207;
  assign T207 = ~ maskHihgerReq_11;
  assign T208 = noReqMasked & grantUnMasked_11;
  assign grantUnMasked_11 = T209;
  assign T209 = requestVec_11 & T210;
  assign T210 = ~ unMaskHigherReq_11;
  assign io_grant_12 = grant_12;
  assign grant_12 = T211;
  assign T211 = T214 | grantMasked_12;
  assign grantMasked_12 = T212;
  assign T212 = requestMasked_12 & T213;
  assign T213 = ~ maskHihgerReq_12;
  assign T214 = noReqMasked & grantUnMasked_12;
  assign grantUnMasked_12 = T215;
  assign T215 = requestVec_12 & T216;
  assign T216 = ~ unMaskHigherReq_12;
  assign io_grant_13 = grant_13;
  assign grant_13 = T217;
  assign T217 = T220 | grantMasked_13;
  assign grantMasked_13 = T218;
  assign T218 = requestMasked_13 & T219;
  assign T219 = ~ maskHihgerReq_13;
  assign T220 = noReqMasked & grantUnMasked_13;
  assign grantUnMasked_13 = T221;
  assign T221 = requestVec_13 & T222;
  assign T222 = ~ unMaskHigherReq_13;
  assign io_grant_14 = grant_14;
  assign grant_14 = T223;
  assign T223 = T226 | grantMasked_14;
  assign grantMasked_14 = T224;
  assign T224 = requestMasked_14 & T225;
  assign T225 = ~ maskHihgerReq_14;
  assign T226 = noReqMasked & grantUnMasked_14;
  assign grantUnMasked_14 = T227;
  assign T227 = requestVec_14 & T228;
  assign T228 = ~ unMaskHigherReq_14;
  assign io_grant_15 = grant_15;
  assign grant_15 = T229;
  assign T229 = T232 | grantMasked_15;
  assign grantMasked_15 = T230;
  assign T230 = requestMasked_15 & T231;
  assign T231 = ~ maskHihgerReq_15;
  assign T232 = noReqMasked & grantUnMasked_15;
  assign grantUnMasked_15 = T233;
  assign T233 = requestVec_15 & T234;
  assign T234 = ~ unMaskHigherReq_15;
  assign io_grant_16 = grant_16;
  assign grant_16 = T235;
  assign T235 = T238 | grantMasked_16;
  assign grantMasked_16 = T236;
  assign T236 = requestMasked_16 & T237;
  assign T237 = ~ maskHihgerReq_16;
  assign T238 = noReqMasked & grantUnMasked_16;
  assign grantUnMasked_16 = T239;
  assign T239 = requestVec_16 & T240;
  assign T240 = ~ unMaskHigherReq_16;
  assign io_grant_17 = grant_17;
  assign grant_17 = T241;
  assign T241 = T244 | grantMasked_17;
  assign grantMasked_17 = T242;
  assign T242 = requestMasked_17 & T243;
  assign T243 = ~ maskHihgerReq_17;
  assign T244 = noReqMasked & grantUnMasked_17;
  assign grantUnMasked_17 = T245;
  assign T245 = requestVec_17 & T246;
  assign T246 = ~ unMaskHigherReq_17;
  assign io_grant_18 = grant_18;
  assign grant_18 = T247;
  assign T247 = T250 | grantMasked_18;
  assign grantMasked_18 = T248;
  assign T248 = requestMasked_18 & T249;
  assign T249 = ~ maskHihgerReq_18;
  assign T250 = noReqMasked & grantUnMasked_18;
  assign grantUnMasked_18 = T251;
  assign T251 = requestVec_18 & T252;
  assign T252 = ~ unMaskHigherReq_18;
  assign io_grant_19 = grant_19;
  assign grant_19 = T253;
  assign T253 = T256 | grantMasked_19;
  assign grantMasked_19 = T254;
  assign T254 = requestMasked_19 & T255;
  assign T255 = ~ maskHihgerReq_19;
  assign T256 = noReqMasked & grantUnMasked_19;
  assign grantUnMasked_19 = T257;
  assign T257 = requestVec_19 & T258;
  assign T258 = ~ unMaskHigherReq_19;

  always @(posedge clk) begin
    if(reset) begin
      pointerReg_0 <= 1'h0;
    end else if(T120) begin
      pointerReg_0 <= unMaskHigherReq_0;
    end else if(anyReqMasked) begin
      pointerReg_0 <= maskHihgerReq_0;
    end
    if(reset) begin
      pointerReg_19 <= 1'h0;
    end else if(T120) begin
      pointerReg_19 <= unMaskHigherReq_19;
    end else if(anyReqMasked) begin
      pointerReg_19 <= maskHihgerReq_19;
    end
    if(reset) begin
      pointerReg_18 <= 1'h0;
    end else if(T120) begin
      pointerReg_18 <= unMaskHigherReq_18;
    end else if(anyReqMasked) begin
      pointerReg_18 <= maskHihgerReq_18;
    end
    if(reset) begin
      pointerReg_17 <= 1'h0;
    end else if(T120) begin
      pointerReg_17 <= unMaskHigherReq_17;
    end else if(anyReqMasked) begin
      pointerReg_17 <= maskHihgerReq_17;
    end
    if(reset) begin
      pointerReg_16 <= 1'h0;
    end else if(T120) begin
      pointerReg_16 <= unMaskHigherReq_16;
    end else if(anyReqMasked) begin
      pointerReg_16 <= maskHihgerReq_16;
    end
    if(reset) begin
      pointerReg_15 <= 1'h0;
    end else if(T120) begin
      pointerReg_15 <= unMaskHigherReq_15;
    end else if(anyReqMasked) begin
      pointerReg_15 <= maskHihgerReq_15;
    end
    if(reset) begin
      pointerReg_14 <= 1'h0;
    end else if(T120) begin
      pointerReg_14 <= unMaskHigherReq_14;
    end else if(anyReqMasked) begin
      pointerReg_14 <= maskHihgerReq_14;
    end
    if(reset) begin
      pointerReg_13 <= 1'h0;
    end else if(T120) begin
      pointerReg_13 <= unMaskHigherReq_13;
    end else if(anyReqMasked) begin
      pointerReg_13 <= maskHihgerReq_13;
    end
    if(reset) begin
      pointerReg_12 <= 1'h0;
    end else if(T120) begin
      pointerReg_12 <= unMaskHigherReq_12;
    end else if(anyReqMasked) begin
      pointerReg_12 <= maskHihgerReq_12;
    end
    if(reset) begin
      pointerReg_11 <= 1'h0;
    end else if(T120) begin
      pointerReg_11 <= unMaskHigherReq_11;
    end else if(anyReqMasked) begin
      pointerReg_11 <= maskHihgerReq_11;
    end
    if(reset) begin
      pointerReg_10 <= 1'h0;
    end else if(T120) begin
      pointerReg_10 <= unMaskHigherReq_10;
    end else if(anyReqMasked) begin
      pointerReg_10 <= maskHihgerReq_10;
    end
    if(reset) begin
      pointerReg_9 <= 1'h0;
    end else if(T120) begin
      pointerReg_9 <= unMaskHigherReq_9;
    end else if(anyReqMasked) begin
      pointerReg_9 <= maskHihgerReq_9;
    end
    if(reset) begin
      pointerReg_8 <= 1'h0;
    end else if(T120) begin
      pointerReg_8 <= unMaskHigherReq_8;
    end else if(anyReqMasked) begin
      pointerReg_8 <= maskHihgerReq_8;
    end
    if(reset) begin
      pointerReg_7 <= 1'h0;
    end else if(T120) begin
      pointerReg_7 <= unMaskHigherReq_7;
    end else if(anyReqMasked) begin
      pointerReg_7 <= maskHihgerReq_7;
    end
    if(reset) begin
      pointerReg_6 <= 1'h0;
    end else if(T120) begin
      pointerReg_6 <= unMaskHigherReq_6;
    end else if(anyReqMasked) begin
      pointerReg_6 <= maskHihgerReq_6;
    end
    if(reset) begin
      pointerReg_5 <= 1'h0;
    end else if(T120) begin
      pointerReg_5 <= unMaskHigherReq_5;
    end else if(anyReqMasked) begin
      pointerReg_5 <= maskHihgerReq_5;
    end
    if(reset) begin
      pointerReg_4 <= 1'h0;
    end else if(T120) begin
      pointerReg_4 <= unMaskHigherReq_4;
    end else if(anyReqMasked) begin
      pointerReg_4 <= maskHihgerReq_4;
    end
    if(reset) begin
      pointerReg_3 <= 1'h0;
    end else if(T120) begin
      pointerReg_3 <= unMaskHigherReq_3;
    end else if(anyReqMasked) begin
      pointerReg_3 <= maskHihgerReq_3;
    end
    if(reset) begin
      pointerReg_2 <= 1'h0;
    end else if(T120) begin
      pointerReg_2 <= unMaskHigherReq_2;
    end else if(anyReqMasked) begin
      pointerReg_2 <= maskHihgerReq_2;
    end
    if(reset) begin
      pointerReg_1 <= 1'h0;
    end else if(T120) begin
      pointerReg_1 <= unMaskHigherReq_1;
    end else if(anyReqMasked) begin
      pointerReg_1 <= maskHihgerReq_1;
    end
  end
endmodule

module fifoFabOut_0(input clk, input reset,
    input [55:0] io_enqData,
    output[55:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    output[1:0] io_emptySpace,
    input  io_rst
);

  wire[1:0] emptySpace;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire isFullNext;
  wire T7;
  reg  isFull;
  wire T80;
  wire T8;
  wire rst;
  wire T9;
  wire doDeq;
  wire T10;
  wire T11;
  wire T12;
  reg [1:0] deqPtr;
  wire[1:0] T81;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] deqPtrInc;
  wire[1:0] T15;
  wire[1:0] enqPtrInc;
  wire[1:0] T16;
  reg [1:0] enqPtr;
  wire[1:0] T82;
  wire[1:0] T17;
  wire[1:0] T18;
  wire doEnq;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire isEmpty;
  wire T72;
  wire T73;
  wire T74;
  wire[55:0] T75;
  reg [55:0] fifoMem [2:0];
  wire[55:0] T76;
  wire T77;
  wire T78;
  wire[1:0] T79;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    isFull = {1{$random}};
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_emptySpace = emptySpace;
  assign emptySpace = T0;
  assign T0 = T63 ? T62 : T1;
  assign T1 = T54 ? T53 : T2;
  assign T2 = T46 ? T45 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T30 ? T29 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = isFullNext ? 2'h0 : 2'h3;
  assign isFullNext = T11 ? 1'h1 : T7;
  assign T7 = T9 ? 1'h0 : isFull;
  assign T80 = reset ? 1'h0 : T8;
  assign T8 = rst ? 1'h0 : isFullNext;
  assign rst = io_rst;
  assign T9 = doDeq & isFull;
  assign doDeq = T10;
  assign T10 = io_deqValid & io_deqRdy;
  assign T11 = T20 & T12;
  assign T12 = enqPtrInc == deqPtr;
  assign T81 = reset ? 2'h0 : T13;
  assign T13 = rst ? 2'h0 : T14;
  assign T14 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T15 % 2'h3;
  assign T15 = deqPtr + 2'h1;
  assign enqPtrInc = T16 % 2'h3;
  assign T16 = enqPtr + 2'h1;
  assign T82 = reset ? 2'h0 : T17;
  assign T17 = rst ? 2'h0 : T18;
  assign T18 = doEnq ? enqPtrInc : enqPtr;
  assign doEnq = T19;
  assign T19 = io_enqRdy & io_enqValid;
  assign T20 = doEnq & T21;
  assign T21 = ~ doDeq;
  assign T22 = enqPtrInc - deqPtr;
  assign T23 = T28 & T24;
  assign T24 = T26 & T25;
  assign T25 = deqPtr < enqPtrInc;
  assign T26 = doEnq & T27;
  assign T27 = ~ doDeq;
  assign T28 = isFullNext ^ 1'h1;
  assign T29 = deqPtr - enqPtrInc;
  assign T30 = T35 & T31;
  assign T31 = T33 & T32;
  assign T32 = enqPtrInc < deqPtr;
  assign T33 = doEnq & T34;
  assign T34 = ~ doDeq;
  assign T35 = T36 ^ 1'h1;
  assign T36 = isFullNext | T24;
  assign T37 = enqPtr - deqPtrInc;
  assign T38 = T43 & T39;
  assign T39 = T41 & T40;
  assign T40 = deqPtrInc < enqPtr;
  assign T41 = T42 & doDeq;
  assign T42 = ~ doEnq;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T36 | T31;
  assign T45 = deqPtrInc - enqPtr;
  assign T46 = T51 & T47;
  assign T47 = T49 & T48;
  assign T48 = enqPtr < deqPtrInc;
  assign T49 = T50 & doDeq;
  assign T50 = ~ doEnq;
  assign T51 = T52 ^ 1'h1;
  assign T52 = T44 | T39;
  assign T53 = enqPtr - deqPtr;
  assign T54 = T60 & T55;
  assign T55 = T57 & T56;
  assign T56 = deqPtr < enqPtr;
  assign T57 = T59 & T58;
  assign T58 = ~ doDeq;
  assign T59 = ~ doEnq;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T52 | T47;
  assign T62 = deqPtr - enqPtr;
  assign T63 = T69 & T64;
  assign T64 = T66 & T65;
  assign T65 = enqPtr < deqPtr;
  assign T66 = T68 & T67;
  assign T67 = ~ doDeq;
  assign T68 = ~ doEnq;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T61 | T55;
  assign io_deqValid = T71;
  assign T71 = isEmpty ^ 1'h1;
  assign isEmpty = T73 & T72;
  assign T72 = enqPtr == deqPtr;
  assign T73 = isFull ^ 1'h1;
  assign io_enqRdy = T74;
  assign T74 = isFull ^ 1'h1;
  assign io_deqData = T75;
  assign T75 = fifoMem[deqPtr];
  assign T77 = doEnq & T78;
  assign T78 = T79 < 2'h3;
  assign T79 = enqPtr[1'h1:1'h0];

  always @(posedge clk) begin
    if(reset) begin
      isFull <= 1'h0;
    end else if(rst) begin
      isFull <= 1'h0;
    end else if(T11) begin
      isFull <= 1'h1;
    end else if(T9) begin
      isFull <= 1'h0;
    end
    if(reset) begin
      deqPtr <= 2'h0;
    end else if(rst) begin
      deqPtr <= 2'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 2'h0;
    end else if(rst) begin
      enqPtr <= 2'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if (T77)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fifoFabOut_1(input clk, input reset,
    input [55:0] io_enqData,
    output[55:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    output[1:0] io_emptySpace,
    input  io_rst
);

  wire[1:0] emptySpace;
  wire[1:0] T77;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire isFullNext;
  wire T7;
  reg  isFull;
  wire T78;
  wire T8;
  wire rst;
  wire T9;
  wire doDeq;
  wire T10;
  wire T11;
  wire T12;
  reg [1:0] deqPtr;
  wire[1:0] T79;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] deqPtrInc;
  wire[1:0] T15;
  wire[1:0] enqPtrInc;
  wire[1:0] T16;
  reg [1:0] enqPtr;
  wire[1:0] T80;
  wire[1:0] T17;
  wire[1:0] T18;
  wire doEnq;
  wire T19;
  wire T20;
  wire T21;
  wire[2:0] T81;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[2:0] T82;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[2:0] T83;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[2:0] T84;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[2:0] T85;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T86;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire isEmpty;
  wire T72;
  wire T73;
  wire T74;
  wire[55:0] T75;
  reg [55:0] fifoMem [3:0];
  wire[55:0] T76;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    isFull = {1{$random}};
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_emptySpace = emptySpace;
  assign emptySpace = T77;
  assign T77 = T0[1'h1:1'h0];
  assign T0 = T63 ? T86 : T1;
  assign T1 = T54 ? T85 : T2;
  assign T2 = T46 ? T84 : T3;
  assign T3 = T38 ? T83 : T4;
  assign T4 = T30 ? T82 : T5;
  assign T5 = T23 ? T81 : T6;
  assign T6 = isFullNext ? 3'h0 : 3'h4;
  assign isFullNext = T11 ? 1'h1 : T7;
  assign T7 = T9 ? 1'h0 : isFull;
  assign T78 = reset ? 1'h0 : T8;
  assign T8 = rst ? 1'h0 : isFullNext;
  assign rst = io_rst;
  assign T9 = doDeq & isFull;
  assign doDeq = T10;
  assign T10 = io_deqValid & io_deqRdy;
  assign T11 = T20 & T12;
  assign T12 = enqPtrInc == deqPtr;
  assign T79 = reset ? 2'h0 : T13;
  assign T13 = rst ? 2'h0 : T14;
  assign T14 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T15 % 3'h4;
  assign T15 = deqPtr + 2'h1;
  assign enqPtrInc = T16 % 3'h4;
  assign T16 = enqPtr + 2'h1;
  assign T80 = reset ? 2'h0 : T17;
  assign T17 = rst ? 2'h0 : T18;
  assign T18 = doEnq ? enqPtrInc : enqPtr;
  assign doEnq = T19;
  assign T19 = io_enqRdy & io_enqValid;
  assign T20 = doEnq & T21;
  assign T21 = ~ doDeq;
  assign T81 = {1'h0, T22};
  assign T22 = enqPtrInc - deqPtr;
  assign T23 = T28 & T24;
  assign T24 = T26 & T25;
  assign T25 = deqPtr < enqPtrInc;
  assign T26 = doEnq & T27;
  assign T27 = ~ doDeq;
  assign T28 = isFullNext ^ 1'h1;
  assign T82 = {1'h0, T29};
  assign T29 = deqPtr - enqPtrInc;
  assign T30 = T35 & T31;
  assign T31 = T33 & T32;
  assign T32 = enqPtrInc < deqPtr;
  assign T33 = doEnq & T34;
  assign T34 = ~ doDeq;
  assign T35 = T36 ^ 1'h1;
  assign T36 = isFullNext | T24;
  assign T83 = {1'h0, T37};
  assign T37 = enqPtr - deqPtrInc;
  assign T38 = T43 & T39;
  assign T39 = T41 & T40;
  assign T40 = deqPtrInc < enqPtr;
  assign T41 = T42 & doDeq;
  assign T42 = ~ doEnq;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T36 | T31;
  assign T84 = {1'h0, T45};
  assign T45 = deqPtrInc - enqPtr;
  assign T46 = T51 & T47;
  assign T47 = T49 & T48;
  assign T48 = enqPtr < deqPtrInc;
  assign T49 = T50 & doDeq;
  assign T50 = ~ doEnq;
  assign T51 = T52 ^ 1'h1;
  assign T52 = T44 | T39;
  assign T85 = {1'h0, T53};
  assign T53 = enqPtr - deqPtr;
  assign T54 = T60 & T55;
  assign T55 = T57 & T56;
  assign T56 = deqPtr < enqPtr;
  assign T57 = T59 & T58;
  assign T58 = ~ doDeq;
  assign T59 = ~ doEnq;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T52 | T47;
  assign T86 = {1'h0, T62};
  assign T62 = deqPtr - enqPtr;
  assign T63 = T69 & T64;
  assign T64 = T66 & T65;
  assign T65 = enqPtr < deqPtr;
  assign T66 = T68 & T67;
  assign T67 = ~ doDeq;
  assign T68 = ~ doEnq;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T61 | T55;
  assign io_deqValid = T71;
  assign T71 = isEmpty ^ 1'h1;
  assign isEmpty = T73 & T72;
  assign T72 = enqPtr == deqPtr;
  assign T73 = isFull ^ 1'h1;
  assign io_enqRdy = T74;
  assign T74 = isFull ^ 1'h1;
  assign io_deqData = T75;
  assign T75 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      isFull <= 1'h0;
    end else if(rst) begin
      isFull <= 1'h0;
    end else if(T11) begin
      isFull <= 1'h1;
    end else if(T9) begin
      isFull <= 1'h0;
    end
    if(reset) begin
      deqPtr <= 2'h0;
    end else if(rst) begin
      deqPtr <= 2'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 2'h0;
    end else if(rst) begin
      enqPtr <= 2'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fabOutSeqArb(input clk, input reset,
    input [55:0] io_fabOutLoc_19,
    input [55:0] io_fabOutLoc_18,
    input [55:0] io_fabOutLoc_17,
    input [55:0] io_fabOutLoc_16,
    input [55:0] io_fabOutLoc_15,
    input [55:0] io_fabOutLoc_14,
    input [55:0] io_fabOutLoc_13,
    input [55:0] io_fabOutLoc_12,
    input [55:0] io_fabOutLoc_11,
    input [55:0] io_fabOutLoc_10,
    input [55:0] io_fabOutLoc_9,
    input [55:0] io_fabOutLoc_8,
    input [55:0] io_fabOutLoc_7,
    input [55:0] io_fabOutLoc_6,
    input [55:0] io_fabOutLoc_5,
    input [55:0] io_fabOutLoc_4,
    input [55:0] io_fabOutLoc_3,
    input [55:0] io_fabOutLoc_2,
    input [55:0] io_fabOutLoc_1,
    input [55:0] io_fabOutLoc_0,
    input  io_fabOutLocValid_19,
    input  io_fabOutLocValid_18,
    input  io_fabOutLocValid_17,
    input  io_fabOutLocValid_16,
    input  io_fabOutLocValid_15,
    input  io_fabOutLocValid_14,
    input  io_fabOutLocValid_13,
    input  io_fabOutLocValid_12,
    input  io_fabOutLocValid_11,
    input  io_fabOutLocValid_10,
    input  io_fabOutLocValid_9,
    input  io_fabOutLocValid_8,
    input  io_fabOutLocValid_7,
    input  io_fabOutLocValid_6,
    input  io_fabOutLocValid_5,
    input  io_fabOutLocValid_4,
    input  io_fabOutLocValid_3,
    input  io_fabOutLocValid_2,
    input  io_fabOutLocValid_1,
    input  io_fabOutLocValid_0,
    output io_fabOutLocRdy_19,
    output io_fabOutLocRdy_18,
    output io_fabOutLocRdy_17,
    output io_fabOutLocRdy_16,
    output io_fabOutLocRdy_15,
    output io_fabOutLocRdy_14,
    output io_fabOutLocRdy_13,
    output io_fabOutLocRdy_12,
    output io_fabOutLocRdy_11,
    output io_fabOutLocRdy_10,
    output io_fabOutLocRdy_9,
    output io_fabOutLocRdy_8,
    output io_fabOutLocRdy_7,
    output io_fabOutLocRdy_6,
    output io_fabOutLocRdy_5,
    output io_fabOutLocRdy_4,
    output io_fabOutLocRdy_3,
    output io_fabOutLocRdy_2,
    output io_fabOutLocRdy_1,
    output io_fabOutLocRdy_0,
    output[55:0] io_locStoreData,
    output io_locStoreValid,
    input  io_locStoreRdy,
    input  io_rst
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg  muxValidReg_0;
  wire T341;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg  grantReg_0;
  wire T342;
  wire grantWire_0;
  reg  grantReg_1;
  wire T343;
  wire grantWire_1;
  reg  grantReg_2;
  wire T344;
  wire grantWire_2;
  reg  grantReg_3;
  wire T345;
  wire grantWire_3;
  wire T19;
  reg  muxValidReg_1;
  wire T346;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  grantReg_4;
  wire T347;
  wire grantWire_4;
  reg  grantReg_5;
  wire T348;
  wire grantWire_5;
  reg  grantReg_6;
  wire T349;
  wire grantWire_6;
  reg  grantReg_7;
  wire T350;
  wire grantWire_7;
  wire T29;
  wire T30;
  reg  muxValidReg_2;
  wire T351;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg  grantReg_8;
  wire T352;
  wire grantWire_8;
  reg  grantReg_9;
  wire T353;
  wire grantWire_9;
  reg  grantReg_10;
  wire T354;
  wire grantWire_10;
  reg  grantReg_11;
  wire T355;
  wire grantWire_11;
  wire T40;
  wire T41;
  reg  muxValidReg_3;
  wire T356;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  grantReg_12;
  wire T357;
  wire grantWire_12;
  reg  grantReg_13;
  wire T358;
  wire grantWire_13;
  reg  grantReg_14;
  wire T359;
  wire grantWire_14;
  reg  grantReg_15;
  wire T360;
  wire grantWire_15;
  wire T51;
  wire T52;
  reg  muxValidReg_4;
  wire T361;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  reg  grantReg_16;
  wire T362;
  wire grantWire_16;
  reg  grantReg_17;
  wire T363;
  wire grantWire_17;
  reg  grantReg_18;
  wire T364;
  wire grantWire_18;
  reg  grantReg_19;
  wire T365;
  wire grantWire_19;
  wire T62;
  wire T63;
  wire[55:0] T64;
  wire[55:0] T65;
  wire[55:0] T66;
  wire[55:0] T67;
  wire[55:0] T68;
  wire[55:0] T69;
  wire[55:0] T70;
  wire[55:0] T71;
  wire[55:0] T72;
  reg [55:0] muxReg_0;
  wire[55:0] T366;
  wire[55:0] T73;
  wire[55:0] T74;
  wire[55:0] T75;
  wire[55:0] T76;
  reg [55:0] muxReg_1;
  wire[55:0] T367;
  wire[55:0] T77;
  wire[55:0] T78;
  wire[55:0] T79;
  wire[55:0] T80;
  reg [55:0] muxReg_2;
  wire[55:0] T368;
  wire[55:0] T81;
  wire[55:0] T82;
  wire[55:0] T83;
  wire[55:0] T84;
  reg [55:0] muxReg_3;
  wire[55:0] T369;
  wire[55:0] T85;
  wire[55:0] T86;
  wire[55:0] T87;
  wire[55:0] T88;
  reg [55:0] muxReg_4;
  wire[55:0] T370;
  wire[55:0] T89;
  wire[55:0] T90;
  wire[55:0] T91;
  wire[55:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire request_0;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire anyGrant;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire muxValid;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire request_1;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire request_2;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire request_3;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire request_4;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire request_5;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire request_6;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire request_7;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire request_8;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire request_9;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire request_10;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire request_11;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire request_12;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire request_13;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire request_14;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire request_15;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire request_16;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire request_17;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire request_18;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire request_19;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire arb_io_grant_19;
  wire arb_io_grant_18;
  wire arb_io_grant_17;
  wire arb_io_grant_16;
  wire arb_io_grant_15;
  wire arb_io_grant_14;
  wire arb_io_grant_13;
  wire arb_io_grant_12;
  wire arb_io_grant_11;
  wire arb_io_grant_10;
  wire arb_io_grant_9;
  wire arb_io_grant_8;
  wire arb_io_grant_7;
  wire arb_io_grant_6;
  wire arb_io_grant_5;
  wire arb_io_grant_4;
  wire arb_io_grant_3;
  wire arb_io_grant_2;
  wire arb_io_grant_1;
  wire arb_io_grant_0;
  wire[55:0] fifoFabOut_io_deqData;
  wire fifoFabOut_io_enqRdy;
  wire fifoFabOut_io_deqValid;
  wire[1:0] fifoFabOut_io_emptySpace;
  wire[55:0] fifoFabOut_1_io_deqData;
  wire fifoFabOut_1_io_enqRdy;
  wire fifoFabOut_1_io_deqValid;
  wire[1:0] fifoFabOut_1_io_emptySpace;
  wire[55:0] fifoFabOut_2_io_deqData;
  wire fifoFabOut_2_io_enqRdy;
  wire fifoFabOut_2_io_deqValid;
  wire[1:0] fifoFabOut_2_io_emptySpace;
  wire[55:0] fifoFabOut_3_io_deqData;
  wire fifoFabOut_3_io_enqRdy;
  wire fifoFabOut_3_io_deqValid;
  wire[1:0] fifoFabOut_3_io_emptySpace;
  wire[55:0] fifoFabOut_4_io_deqData;
  wire fifoFabOut_4_io_enqRdy;
  wire fifoFabOut_4_io_deqValid;
  wire[1:0] fifoFabOut_4_io_emptySpace;
  wire[55:0] fifoFabOut_5_io_deqData;
  wire fifoFabOut_5_io_enqRdy;
  wire fifoFabOut_5_io_deqValid;
  wire[1:0] fifoFabOut_5_io_emptySpace;
  wire[55:0] fifoFabOut_6_io_deqData;
  wire fifoFabOut_6_io_enqRdy;
  wire fifoFabOut_6_io_deqValid;
  wire[1:0] fifoFabOut_6_io_emptySpace;
  wire[55:0] fifoFabOut_7_io_deqData;
  wire fifoFabOut_7_io_enqRdy;
  wire fifoFabOut_7_io_deqValid;
  wire[1:0] fifoFabOut_7_io_emptySpace;
  wire[55:0] fifoFabOut_8_io_deqData;
  wire fifoFabOut_8_io_enqRdy;
  wire fifoFabOut_8_io_deqValid;
  wire[1:0] fifoFabOut_8_io_emptySpace;
  wire[55:0] fifoFabOut_9_io_deqData;
  wire fifoFabOut_9_io_enqRdy;
  wire fifoFabOut_9_io_deqValid;
  wire[1:0] fifoFabOut_9_io_emptySpace;
  wire[55:0] fifoFabOut_10_io_deqData;
  wire fifoFabOut_10_io_enqRdy;
  wire fifoFabOut_10_io_deqValid;
  wire[1:0] fifoFabOut_10_io_emptySpace;
  wire[55:0] fifoFabOut_11_io_deqData;
  wire fifoFabOut_11_io_enqRdy;
  wire fifoFabOut_11_io_deqValid;
  wire[1:0] fifoFabOut_11_io_emptySpace;
  wire[55:0] fifoFabOut_12_io_deqData;
  wire fifoFabOut_12_io_enqRdy;
  wire fifoFabOut_12_io_deqValid;
  wire[1:0] fifoFabOut_12_io_emptySpace;
  wire[55:0] fifoFabOut_13_io_deqData;
  wire fifoFabOut_13_io_enqRdy;
  wire fifoFabOut_13_io_deqValid;
  wire[1:0] fifoFabOut_13_io_emptySpace;
  wire[55:0] fifoFabOut_14_io_deqData;
  wire fifoFabOut_14_io_enqRdy;
  wire fifoFabOut_14_io_deqValid;
  wire[1:0] fifoFabOut_14_io_emptySpace;
  wire[55:0] fifoFabOut_15_io_deqData;
  wire fifoFabOut_15_io_enqRdy;
  wire fifoFabOut_15_io_deqValid;
  wire[1:0] fifoFabOut_15_io_emptySpace;
  wire[55:0] fifoFabOut_16_io_deqData;
  wire fifoFabOut_16_io_enqRdy;
  wire fifoFabOut_16_io_deqValid;
  wire[1:0] fifoFabOut_16_io_emptySpace;
  wire[55:0] fifoFabOut_17_io_deqData;
  wire fifoFabOut_17_io_enqRdy;
  wire fifoFabOut_17_io_deqValid;
  wire[1:0] fifoFabOut_17_io_emptySpace;
  wire[55:0] fifoFabOut_18_io_deqData;
  wire fifoFabOut_18_io_enqRdy;
  wire fifoFabOut_18_io_deqValid;
  wire[1:0] fifoFabOut_18_io_emptySpace;
  wire[55:0] fifoFabOut_19_io_deqData;
  wire fifoFabOut_19_io_enqRdy;
  wire fifoFabOut_19_io_deqValid;
  wire[1:0] fifoFabOut_19_io_emptySpace;
  wire[55:0] outFifo_io_deqData;
  wire outFifo_io_enqRdy;
  wire outFifo_io_deqValid;
  wire[1:0] outFifo_io_emptySpace;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    muxValidReg_0 = {1{$random}};
    grantReg_0 = {1{$random}};
    grantReg_1 = {1{$random}};
    grantReg_2 = {1{$random}};
    grantReg_3 = {1{$random}};
    muxValidReg_1 = {1{$random}};
    grantReg_4 = {1{$random}};
    grantReg_5 = {1{$random}};
    grantReg_6 = {1{$random}};
    grantReg_7 = {1{$random}};
    muxValidReg_2 = {1{$random}};
    grantReg_8 = {1{$random}};
    grantReg_9 = {1{$random}};
    grantReg_10 = {1{$random}};
    grantReg_11 = {1{$random}};
    muxValidReg_3 = {1{$random}};
    grantReg_12 = {1{$random}};
    grantReg_13 = {1{$random}};
    grantReg_14 = {1{$random}};
    grantReg_15 = {1{$random}};
    muxValidReg_4 = {1{$random}};
    grantReg_16 = {1{$random}};
    grantReg_17 = {1{$random}};
    grantReg_18 = {1{$random}};
    grantReg_19 = {1{$random}};
    muxReg_0 = {2{$random}};
    muxReg_1 = {2{$random}};
    muxReg_2 = {2{$random}};
    muxReg_3 = {2{$random}};
    muxReg_4 = {2{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_rst ? 1'h1 : 1'h0;
  assign T1 = T63 ? 1'h0 : T2;
  assign T2 = T62 ? muxValidReg_4 : T3;
  assign T3 = T52 ? 1'h0 : T4;
  assign T4 = T51 ? muxValidReg_3 : T5;
  assign T5 = T41 ? 1'h0 : T6;
  assign T6 = T40 ? muxValidReg_2 : T7;
  assign T7 = T30 ? 1'h0 : T8;
  assign T8 = T29 ? muxValidReg_1 : T9;
  assign T9 = T19 ? muxValidReg_0 : 1'h0;
  assign T341 = reset ? 1'h0 : T10;
  assign T10 = io_rst ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : T12;
  assign T12 = io_rst ? 1'h0 : T13;
  assign T13 = io_rst ? 1'h0 : T14;
  assign T14 = io_rst ? 1'h0 : T15;
  assign T15 = grantReg_3 ? fifoFabOut_3_io_deqValid : T16;
  assign T16 = grantReg_2 ? fifoFabOut_2_io_deqValid : T17;
  assign T17 = grantReg_1 ? fifoFabOut_1_io_deqValid : T18;
  assign T18 = grantReg_0 ? fifoFabOut_io_deqValid : muxValidReg_0;
  assign T342 = reset ? 1'h0 : grantWire_0;
  assign grantWire_0 = arb_io_grant_0;
  assign T343 = reset ? 1'h0 : grantWire_1;
  assign grantWire_1 = arb_io_grant_1;
  assign T344 = reset ? 1'h0 : grantWire_2;
  assign grantWire_2 = arb_io_grant_2;
  assign T345 = reset ? 1'h0 : grantWire_3;
  assign grantWire_3 = arb_io_grant_3;
  assign T19 = muxValidReg_0 & outFifo_io_enqRdy;
  assign T346 = reset ? 1'h0 : T20;
  assign T20 = io_rst ? 1'h0 : T21;
  assign T21 = io_rst ? 1'h0 : T22;
  assign T22 = io_rst ? 1'h0 : T23;
  assign T23 = io_rst ? 1'h0 : T24;
  assign T24 = io_rst ? 1'h0 : T25;
  assign T25 = grantReg_7 ? fifoFabOut_7_io_deqValid : T26;
  assign T26 = grantReg_6 ? fifoFabOut_6_io_deqValid : T27;
  assign T27 = grantReg_5 ? fifoFabOut_5_io_deqValid : T28;
  assign T28 = grantReg_4 ? fifoFabOut_4_io_deqValid : muxValidReg_1;
  assign T347 = reset ? 1'h0 : grantWire_4;
  assign grantWire_4 = arb_io_grant_4;
  assign T348 = reset ? 1'h0 : grantWire_5;
  assign grantWire_5 = arb_io_grant_5;
  assign T349 = reset ? 1'h0 : grantWire_6;
  assign grantWire_6 = arb_io_grant_6;
  assign T350 = reset ? 1'h0 : grantWire_7;
  assign grantWire_7 = arb_io_grant_7;
  assign T29 = muxValidReg_1 & outFifo_io_enqRdy;
  assign T30 = T29 ^ 1'h1;
  assign T351 = reset ? 1'h0 : T31;
  assign T31 = io_rst ? 1'h0 : T32;
  assign T32 = io_rst ? 1'h0 : T33;
  assign T33 = io_rst ? 1'h0 : T34;
  assign T34 = io_rst ? 1'h0 : T35;
  assign T35 = io_rst ? 1'h0 : T36;
  assign T36 = grantReg_11 ? fifoFabOut_11_io_deqValid : T37;
  assign T37 = grantReg_10 ? fifoFabOut_10_io_deqValid : T38;
  assign T38 = grantReg_9 ? fifoFabOut_9_io_deqValid : T39;
  assign T39 = grantReg_8 ? fifoFabOut_8_io_deqValid : muxValidReg_2;
  assign T352 = reset ? 1'h0 : grantWire_8;
  assign grantWire_8 = arb_io_grant_8;
  assign T353 = reset ? 1'h0 : grantWire_9;
  assign grantWire_9 = arb_io_grant_9;
  assign T354 = reset ? 1'h0 : grantWire_10;
  assign grantWire_10 = arb_io_grant_10;
  assign T355 = reset ? 1'h0 : grantWire_11;
  assign grantWire_11 = arb_io_grant_11;
  assign T40 = muxValidReg_2 & outFifo_io_enqRdy;
  assign T41 = T40 ^ 1'h1;
  assign T356 = reset ? 1'h0 : T42;
  assign T42 = io_rst ? 1'h0 : T43;
  assign T43 = io_rst ? 1'h0 : T44;
  assign T44 = io_rst ? 1'h0 : T45;
  assign T45 = io_rst ? 1'h0 : T46;
  assign T46 = io_rst ? 1'h0 : T47;
  assign T47 = grantReg_15 ? fifoFabOut_15_io_deqValid : T48;
  assign T48 = grantReg_14 ? fifoFabOut_14_io_deqValid : T49;
  assign T49 = grantReg_13 ? fifoFabOut_13_io_deqValid : T50;
  assign T50 = grantReg_12 ? fifoFabOut_12_io_deqValid : muxValidReg_3;
  assign T357 = reset ? 1'h0 : grantWire_12;
  assign grantWire_12 = arb_io_grant_12;
  assign T358 = reset ? 1'h0 : grantWire_13;
  assign grantWire_13 = arb_io_grant_13;
  assign T359 = reset ? 1'h0 : grantWire_14;
  assign grantWire_14 = arb_io_grant_14;
  assign T360 = reset ? 1'h0 : grantWire_15;
  assign grantWire_15 = arb_io_grant_15;
  assign T51 = muxValidReg_3 & outFifo_io_enqRdy;
  assign T52 = T51 ^ 1'h1;
  assign T361 = reset ? 1'h0 : T53;
  assign T53 = io_rst ? 1'h0 : T54;
  assign T54 = io_rst ? 1'h0 : T55;
  assign T55 = io_rst ? 1'h0 : T56;
  assign T56 = io_rst ? 1'h0 : T57;
  assign T57 = io_rst ? 1'h0 : T58;
  assign T58 = grantReg_19 ? fifoFabOut_19_io_deqValid : T59;
  assign T59 = grantReg_18 ? fifoFabOut_18_io_deqValid : T60;
  assign T60 = grantReg_17 ? fifoFabOut_17_io_deqValid : T61;
  assign T61 = grantReg_16 ? fifoFabOut_16_io_deqValid : muxValidReg_4;
  assign T362 = reset ? 1'h0 : grantWire_16;
  assign grantWire_16 = arb_io_grant_16;
  assign T363 = reset ? 1'h0 : grantWire_17;
  assign grantWire_17 = arb_io_grant_17;
  assign T364 = reset ? 1'h0 : grantWire_18;
  assign grantWire_18 = arb_io_grant_18;
  assign T365 = reset ? 1'h0 : grantWire_19;
  assign grantWire_19 = arb_io_grant_19;
  assign T62 = muxValidReg_4 & outFifo_io_enqRdy;
  assign T63 = T62 ^ 1'h1;
  assign T64 = T63 ? muxReg_4 : T65;
  assign T65 = T62 ? muxReg_4 : T66;
  assign T66 = T52 ? muxReg_3 : T67;
  assign T67 = T51 ? muxReg_3 : T68;
  assign T68 = T41 ? muxReg_2 : T69;
  assign T69 = T40 ? muxReg_2 : T70;
  assign T70 = T30 ? muxReg_1 : T71;
  assign T71 = T29 ? muxReg_1 : T72;
  assign T72 = T19 ? muxReg_0 : muxReg_0;
  assign T366 = reset ? 56'h0 : T73;
  assign T73 = grantReg_3 ? fifoFabOut_3_io_deqData : T74;
  assign T74 = grantReg_2 ? fifoFabOut_2_io_deqData : T75;
  assign T75 = grantReg_1 ? fifoFabOut_1_io_deqData : T76;
  assign T76 = grantReg_0 ? fifoFabOut_io_deqData : muxReg_0;
  assign T367 = reset ? 56'h0 : T77;
  assign T77 = grantReg_7 ? fifoFabOut_7_io_deqData : T78;
  assign T78 = grantReg_6 ? fifoFabOut_6_io_deqData : T79;
  assign T79 = grantReg_5 ? fifoFabOut_5_io_deqData : T80;
  assign T80 = grantReg_4 ? fifoFabOut_4_io_deqData : muxReg_1;
  assign T368 = reset ? 56'h0 : T81;
  assign T81 = grantReg_11 ? fifoFabOut_11_io_deqData : T82;
  assign T82 = grantReg_10 ? fifoFabOut_10_io_deqData : T83;
  assign T83 = grantReg_9 ? fifoFabOut_9_io_deqData : T84;
  assign T84 = grantReg_8 ? fifoFabOut_8_io_deqData : muxReg_2;
  assign T369 = reset ? 56'h0 : T85;
  assign T85 = grantReg_15 ? fifoFabOut_15_io_deqData : T86;
  assign T86 = grantReg_14 ? fifoFabOut_14_io_deqData : T87;
  assign T87 = grantReg_13 ? fifoFabOut_13_io_deqData : T88;
  assign T88 = grantReg_12 ? fifoFabOut_12_io_deqData : muxReg_3;
  assign T370 = reset ? 56'h0 : T89;
  assign T89 = grantReg_19 ? fifoFabOut_19_io_deqData : T90;
  assign T90 = grantReg_18 ? fifoFabOut_18_io_deqData : T91;
  assign T91 = grantReg_17 ? fifoFabOut_17_io_deqData : T92;
  assign T92 = grantReg_16 ? fifoFabOut_16_io_deqData : muxReg_4;
  assign T93 = io_rst ? 1'h1 : 1'h0;
  assign T94 = grantReg_19 ? 1'h1 : 1'h0;
  assign T95 = io_rst ? 1'h1 : 1'h0;
  assign T96 = grantReg_18 ? 1'h1 : 1'h0;
  assign T97 = io_rst ? 1'h1 : 1'h0;
  assign T98 = grantReg_17 ? 1'h1 : 1'h0;
  assign T99 = io_rst ? 1'h1 : 1'h0;
  assign T100 = grantReg_16 ? 1'h1 : 1'h0;
  assign T101 = io_rst ? 1'h1 : 1'h0;
  assign T102 = grantReg_15 ? 1'h1 : 1'h0;
  assign T103 = io_rst ? 1'h1 : 1'h0;
  assign T104 = grantReg_14 ? 1'h1 : 1'h0;
  assign T105 = io_rst ? 1'h1 : 1'h0;
  assign T106 = grantReg_13 ? 1'h1 : 1'h0;
  assign T107 = io_rst ? 1'h1 : 1'h0;
  assign T108 = grantReg_12 ? 1'h1 : 1'h0;
  assign T109 = io_rst ? 1'h1 : 1'h0;
  assign T110 = grantReg_11 ? 1'h1 : 1'h0;
  assign T111 = io_rst ? 1'h1 : 1'h0;
  assign T112 = grantReg_10 ? 1'h1 : 1'h0;
  assign T113 = io_rst ? 1'h1 : 1'h0;
  assign T114 = grantReg_9 ? 1'h1 : 1'h0;
  assign T115 = io_rst ? 1'h1 : 1'h0;
  assign T116 = grantReg_8 ? 1'h1 : 1'h0;
  assign T117 = io_rst ? 1'h1 : 1'h0;
  assign T118 = grantReg_7 ? 1'h1 : 1'h0;
  assign T119 = io_rst ? 1'h1 : 1'h0;
  assign T120 = grantReg_6 ? 1'h1 : 1'h0;
  assign T121 = io_rst ? 1'h1 : 1'h0;
  assign T122 = grantReg_5 ? 1'h1 : 1'h0;
  assign T123 = io_rst ? 1'h1 : 1'h0;
  assign T124 = grantReg_4 ? 1'h1 : 1'h0;
  assign T125 = io_rst ? 1'h1 : 1'h0;
  assign T126 = grantReg_3 ? 1'h1 : 1'h0;
  assign T127 = io_rst ? 1'h1 : 1'h0;
  assign T128 = grantReg_2 ? 1'h1 : 1'h0;
  assign T129 = io_rst ? 1'h1 : 1'h0;
  assign T130 = grantReg_1 ? 1'h1 : 1'h0;
  assign T131 = io_rst ? 1'h1 : 1'h0;
  assign T132 = grantReg_0 ? 1'h1 : 1'h0;
  assign request_0 = T133;
  assign T133 = T168 ? 1'h0 : T134;
  assign T134 = T135 ? 1'h1 : 1'h0;
  assign T135 = T140 & T136;
  assign T136 = fifoFabOut_io_deqValid & T137;
  assign T137 = T138 ^ 1'h1;
  assign T138 = T139 & grantReg_0;
  assign T139 = 2'h1 <= fifoFabOut_io_emptySpace;
  assign T140 = T167 | T141;
  assign T141 = T162 & T142;
  assign T142 = anyGrant ^ 1'h1;
  assign anyGrant = T143;
  assign T143 = T144 | grantReg_19;
  assign T144 = T145 | grantReg_18;
  assign T145 = T146 | grantReg_17;
  assign T146 = T147 | grantReg_16;
  assign T147 = T148 | grantReg_15;
  assign T148 = T149 | grantReg_14;
  assign T149 = T150 | grantReg_13;
  assign T150 = T151 | grantReg_12;
  assign T151 = T152 | grantReg_11;
  assign T152 = T153 | grantReg_10;
  assign T153 = T154 | grantReg_9;
  assign T154 = T155 | grantReg_8;
  assign T155 = T156 | grantReg_7;
  assign T156 = T157 | grantReg_6;
  assign T157 = T158 | grantReg_5;
  assign T158 = T159 | grantReg_4;
  assign T159 = T160 | grantReg_3;
  assign T160 = T161 | grantReg_2;
  assign T161 = grantReg_0 | grantReg_1;
  assign T162 = muxValid ^ 1'h1;
  assign muxValid = T163;
  assign T163 = T164 | muxValidReg_4;
  assign T164 = T165 | muxValidReg_3;
  assign T165 = T166 | muxValidReg_2;
  assign T166 = muxValidReg_0 | muxValidReg_1;
  assign T167 = 2'h1 <= outFifo_io_emptySpace;
  assign T168 = T140 & T169;
  assign T169 = T136 ^ 1'h1;
  assign request_1 = T170;
  assign T170 = T177 ? 1'h0 : T171;
  assign T171 = T172 ? 1'h1 : 1'h0;
  assign T172 = T140 & T173;
  assign T173 = fifoFabOut_1_io_deqValid & T174;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T176 & grantReg_1;
  assign T176 = 2'h1 <= fifoFabOut_1_io_emptySpace;
  assign T177 = T140 & T178;
  assign T178 = T173 ^ 1'h1;
  assign request_2 = T179;
  assign T179 = T186 ? 1'h0 : T180;
  assign T180 = T181 ? 1'h1 : 1'h0;
  assign T181 = T140 & T182;
  assign T182 = fifoFabOut_2_io_deqValid & T183;
  assign T183 = T184 ^ 1'h1;
  assign T184 = T185 & grantReg_2;
  assign T185 = 2'h1 <= fifoFabOut_2_io_emptySpace;
  assign T186 = T140 & T187;
  assign T187 = T182 ^ 1'h1;
  assign request_3 = T188;
  assign T188 = T195 ? 1'h0 : T189;
  assign T189 = T190 ? 1'h1 : 1'h0;
  assign T190 = T140 & T191;
  assign T191 = fifoFabOut_3_io_deqValid & T192;
  assign T192 = T193 ^ 1'h1;
  assign T193 = T194 & grantReg_3;
  assign T194 = 2'h1 <= fifoFabOut_3_io_emptySpace;
  assign T195 = T140 & T196;
  assign T196 = T191 ^ 1'h1;
  assign request_4 = T197;
  assign T197 = T204 ? 1'h0 : T198;
  assign T198 = T199 ? 1'h1 : 1'h0;
  assign T199 = T140 & T200;
  assign T200 = fifoFabOut_4_io_deqValid & T201;
  assign T201 = T202 ^ 1'h1;
  assign T202 = T203 & grantReg_4;
  assign T203 = 2'h1 <= fifoFabOut_4_io_emptySpace;
  assign T204 = T140 & T205;
  assign T205 = T200 ^ 1'h1;
  assign request_5 = T206;
  assign T206 = T213 ? 1'h0 : T207;
  assign T207 = T208 ? 1'h1 : 1'h0;
  assign T208 = T140 & T209;
  assign T209 = fifoFabOut_5_io_deqValid & T210;
  assign T210 = T211 ^ 1'h1;
  assign T211 = T212 & grantReg_5;
  assign T212 = 2'h1 <= fifoFabOut_5_io_emptySpace;
  assign T213 = T140 & T214;
  assign T214 = T209 ^ 1'h1;
  assign request_6 = T215;
  assign T215 = T222 ? 1'h0 : T216;
  assign T216 = T217 ? 1'h1 : 1'h0;
  assign T217 = T140 & T218;
  assign T218 = fifoFabOut_6_io_deqValid & T219;
  assign T219 = T220 ^ 1'h1;
  assign T220 = T221 & grantReg_6;
  assign T221 = 2'h1 <= fifoFabOut_6_io_emptySpace;
  assign T222 = T140 & T223;
  assign T223 = T218 ^ 1'h1;
  assign request_7 = T224;
  assign T224 = T231 ? 1'h0 : T225;
  assign T225 = T226 ? 1'h1 : 1'h0;
  assign T226 = T140 & T227;
  assign T227 = fifoFabOut_7_io_deqValid & T228;
  assign T228 = T229 ^ 1'h1;
  assign T229 = T230 & grantReg_7;
  assign T230 = 2'h1 <= fifoFabOut_7_io_emptySpace;
  assign T231 = T140 & T232;
  assign T232 = T227 ^ 1'h1;
  assign request_8 = T233;
  assign T233 = T240 ? 1'h0 : T234;
  assign T234 = T235 ? 1'h1 : 1'h0;
  assign T235 = T140 & T236;
  assign T236 = fifoFabOut_8_io_deqValid & T237;
  assign T237 = T238 ^ 1'h1;
  assign T238 = T239 & grantReg_8;
  assign T239 = 2'h1 <= fifoFabOut_8_io_emptySpace;
  assign T240 = T140 & T241;
  assign T241 = T236 ^ 1'h1;
  assign request_9 = T242;
  assign T242 = T249 ? 1'h0 : T243;
  assign T243 = T244 ? 1'h1 : 1'h0;
  assign T244 = T140 & T245;
  assign T245 = fifoFabOut_9_io_deqValid & T246;
  assign T246 = T247 ^ 1'h1;
  assign T247 = T248 & grantReg_9;
  assign T248 = 2'h1 <= fifoFabOut_9_io_emptySpace;
  assign T249 = T140 & T250;
  assign T250 = T245 ^ 1'h1;
  assign request_10 = T251;
  assign T251 = T258 ? 1'h0 : T252;
  assign T252 = T253 ? 1'h1 : 1'h0;
  assign T253 = T140 & T254;
  assign T254 = fifoFabOut_10_io_deqValid & T255;
  assign T255 = T256 ^ 1'h1;
  assign T256 = T257 & grantReg_10;
  assign T257 = 2'h1 <= fifoFabOut_10_io_emptySpace;
  assign T258 = T140 & T259;
  assign T259 = T254 ^ 1'h1;
  assign request_11 = T260;
  assign T260 = T267 ? 1'h0 : T261;
  assign T261 = T262 ? 1'h1 : 1'h0;
  assign T262 = T140 & T263;
  assign T263 = fifoFabOut_11_io_deqValid & T264;
  assign T264 = T265 ^ 1'h1;
  assign T265 = T266 & grantReg_11;
  assign T266 = 2'h1 <= fifoFabOut_11_io_emptySpace;
  assign T267 = T140 & T268;
  assign T268 = T263 ^ 1'h1;
  assign request_12 = T269;
  assign T269 = T276 ? 1'h0 : T270;
  assign T270 = T271 ? 1'h1 : 1'h0;
  assign T271 = T140 & T272;
  assign T272 = fifoFabOut_12_io_deqValid & T273;
  assign T273 = T274 ^ 1'h1;
  assign T274 = T275 & grantReg_12;
  assign T275 = 2'h1 <= fifoFabOut_12_io_emptySpace;
  assign T276 = T140 & T277;
  assign T277 = T272 ^ 1'h1;
  assign request_13 = T278;
  assign T278 = T285 ? 1'h0 : T279;
  assign T279 = T280 ? 1'h1 : 1'h0;
  assign T280 = T140 & T281;
  assign T281 = fifoFabOut_13_io_deqValid & T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = T284 & grantReg_13;
  assign T284 = 2'h1 <= fifoFabOut_13_io_emptySpace;
  assign T285 = T140 & T286;
  assign T286 = T281 ^ 1'h1;
  assign request_14 = T287;
  assign T287 = T294 ? 1'h0 : T288;
  assign T288 = T289 ? 1'h1 : 1'h0;
  assign T289 = T140 & T290;
  assign T290 = fifoFabOut_14_io_deqValid & T291;
  assign T291 = T292 ^ 1'h1;
  assign T292 = T293 & grantReg_14;
  assign T293 = 2'h1 <= fifoFabOut_14_io_emptySpace;
  assign T294 = T140 & T295;
  assign T295 = T290 ^ 1'h1;
  assign request_15 = T296;
  assign T296 = T303 ? 1'h0 : T297;
  assign T297 = T298 ? 1'h1 : 1'h0;
  assign T298 = T140 & T299;
  assign T299 = fifoFabOut_15_io_deqValid & T300;
  assign T300 = T301 ^ 1'h1;
  assign T301 = T302 & grantReg_15;
  assign T302 = 2'h1 <= fifoFabOut_15_io_emptySpace;
  assign T303 = T140 & T304;
  assign T304 = T299 ^ 1'h1;
  assign request_16 = T305;
  assign T305 = T312 ? 1'h0 : T306;
  assign T306 = T307 ? 1'h1 : 1'h0;
  assign T307 = T140 & T308;
  assign T308 = fifoFabOut_16_io_deqValid & T309;
  assign T309 = T310 ^ 1'h1;
  assign T310 = T311 & grantReg_16;
  assign T311 = 2'h1 <= fifoFabOut_16_io_emptySpace;
  assign T312 = T140 & T313;
  assign T313 = T308 ^ 1'h1;
  assign request_17 = T314;
  assign T314 = T321 ? 1'h0 : T315;
  assign T315 = T316 ? 1'h1 : 1'h0;
  assign T316 = T140 & T317;
  assign T317 = fifoFabOut_17_io_deqValid & T318;
  assign T318 = T319 ^ 1'h1;
  assign T319 = T320 & grantReg_17;
  assign T320 = 2'h1 <= fifoFabOut_17_io_emptySpace;
  assign T321 = T140 & T322;
  assign T322 = T317 ^ 1'h1;
  assign request_18 = T323;
  assign T323 = T330 ? 1'h0 : T324;
  assign T324 = T325 ? 1'h1 : 1'h0;
  assign T325 = T140 & T326;
  assign T326 = fifoFabOut_18_io_deqValid & T327;
  assign T327 = T328 ^ 1'h1;
  assign T328 = T329 & grantReg_18;
  assign T329 = 2'h1 <= fifoFabOut_18_io_emptySpace;
  assign T330 = T140 & T331;
  assign T331 = T326 ^ 1'h1;
  assign request_19 = T332;
  assign T332 = T339 ? 1'h0 : T333;
  assign T333 = T334 ? 1'h1 : 1'h0;
  assign T334 = T140 & T335;
  assign T335 = fifoFabOut_19_io_deqValid & T336;
  assign T336 = T337 ^ 1'h1;
  assign T337 = T338 & grantReg_19;
  assign T338 = 2'h1 <= fifoFabOut_19_io_emptySpace;
  assign T339 = T140 & T340;
  assign T340 = T335 ^ 1'h1;
  assign io_locStoreValid = outFifo_io_deqValid;
  assign io_locStoreData = outFifo_io_deqData;
  assign io_fabOutLocRdy_0 = fifoFabOut_io_enqRdy;
  assign io_fabOutLocRdy_1 = fifoFabOut_1_io_enqRdy;
  assign io_fabOutLocRdy_2 = fifoFabOut_2_io_enqRdy;
  assign io_fabOutLocRdy_3 = fifoFabOut_3_io_enqRdy;
  assign io_fabOutLocRdy_4 = fifoFabOut_4_io_enqRdy;
  assign io_fabOutLocRdy_5 = fifoFabOut_5_io_enqRdy;
  assign io_fabOutLocRdy_6 = fifoFabOut_6_io_enqRdy;
  assign io_fabOutLocRdy_7 = fifoFabOut_7_io_enqRdy;
  assign io_fabOutLocRdy_8 = fifoFabOut_8_io_enqRdy;
  assign io_fabOutLocRdy_9 = fifoFabOut_9_io_enqRdy;
  assign io_fabOutLocRdy_10 = fifoFabOut_10_io_enqRdy;
  assign io_fabOutLocRdy_11 = fifoFabOut_11_io_enqRdy;
  assign io_fabOutLocRdy_12 = fifoFabOut_12_io_enqRdy;
  assign io_fabOutLocRdy_13 = fifoFabOut_13_io_enqRdy;
  assign io_fabOutLocRdy_14 = fifoFabOut_14_io_enqRdy;
  assign io_fabOutLocRdy_15 = fifoFabOut_15_io_enqRdy;
  assign io_fabOutLocRdy_16 = fifoFabOut_16_io_enqRdy;
  assign io_fabOutLocRdy_17 = fifoFabOut_17_io_enqRdy;
  assign io_fabOutLocRdy_18 = fifoFabOut_18_io_enqRdy;
  assign io_fabOutLocRdy_19 = fifoFabOut_19_io_enqRdy;
  RRArbiter arb(.clk(clk), .reset(reset),
       .io_request_19( request_19 ),
       .io_request_18( request_18 ),
       .io_request_17( request_17 ),
       .io_request_16( request_16 ),
       .io_request_15( request_15 ),
       .io_request_14( request_14 ),
       .io_request_13( request_13 ),
       .io_request_12( request_12 ),
       .io_request_11( request_11 ),
       .io_request_10( request_10 ),
       .io_request_9( request_9 ),
       .io_request_8( request_8 ),
       .io_request_7( request_7 ),
       .io_request_6( request_6 ),
       .io_request_5( request_5 ),
       .io_request_4( request_4 ),
       .io_request_3( request_3 ),
       .io_request_2( request_2 ),
       .io_request_1( request_1 ),
       .io_request_0( request_0 ),
       .io_grant_19( arb_io_grant_19 ),
       .io_grant_18( arb_io_grant_18 ),
       .io_grant_17( arb_io_grant_17 ),
       .io_grant_16( arb_io_grant_16 ),
       .io_grant_15( arb_io_grant_15 ),
       .io_grant_14( arb_io_grant_14 ),
       .io_grant_13( arb_io_grant_13 ),
       .io_grant_12( arb_io_grant_12 ),
       .io_grant_11( arb_io_grant_11 ),
       .io_grant_10( arb_io_grant_10 ),
       .io_grant_9( arb_io_grant_9 ),
       .io_grant_8( arb_io_grant_8 ),
       .io_grant_7( arb_io_grant_7 ),
       .io_grant_6( arb_io_grant_6 ),
       .io_grant_5( arb_io_grant_5 ),
       .io_grant_4( arb_io_grant_4 ),
       .io_grant_3( arb_io_grant_3 ),
       .io_grant_2( arb_io_grant_2 ),
       .io_grant_1( arb_io_grant_1 ),
       .io_grant_0( arb_io_grant_0 )
  );
  fifoFabOut_0 fifoFabOut(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_0 ),
       .io_deqData( fifoFabOut_io_deqData ),
       .io_enqRdy( fifoFabOut_io_enqRdy ),
       .io_deqRdy( T132 ),
       .io_enqValid( io_fabOutLocValid_0 ),
       .io_deqValid( fifoFabOut_io_deqValid ),
       .io_emptySpace( fifoFabOut_io_emptySpace ),
       .io_rst( T131 )
  );
  fifoFabOut_0 fifoFabOut_1(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_1 ),
       .io_deqData( fifoFabOut_1_io_deqData ),
       .io_enqRdy( fifoFabOut_1_io_enqRdy ),
       .io_deqRdy( T130 ),
       .io_enqValid( io_fabOutLocValid_1 ),
       .io_deqValid( fifoFabOut_1_io_deqValid ),
       .io_emptySpace( fifoFabOut_1_io_emptySpace ),
       .io_rst( T129 )
  );
  fifoFabOut_0 fifoFabOut_2(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_2 ),
       .io_deqData( fifoFabOut_2_io_deqData ),
       .io_enqRdy( fifoFabOut_2_io_enqRdy ),
       .io_deqRdy( T128 ),
       .io_enqValid( io_fabOutLocValid_2 ),
       .io_deqValid( fifoFabOut_2_io_deqValid ),
       .io_emptySpace( fifoFabOut_2_io_emptySpace ),
       .io_rst( T127 )
  );
  fifoFabOut_0 fifoFabOut_3(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_3 ),
       .io_deqData( fifoFabOut_3_io_deqData ),
       .io_enqRdy( fifoFabOut_3_io_enqRdy ),
       .io_deqRdy( T126 ),
       .io_enqValid( io_fabOutLocValid_3 ),
       .io_deqValid( fifoFabOut_3_io_deqValid ),
       .io_emptySpace( fifoFabOut_3_io_emptySpace ),
       .io_rst( T125 )
  );
  fifoFabOut_0 fifoFabOut_4(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_4 ),
       .io_deqData( fifoFabOut_4_io_deqData ),
       .io_enqRdy( fifoFabOut_4_io_enqRdy ),
       .io_deqRdy( T124 ),
       .io_enqValid( io_fabOutLocValid_4 ),
       .io_deqValid( fifoFabOut_4_io_deqValid ),
       .io_emptySpace( fifoFabOut_4_io_emptySpace ),
       .io_rst( T123 )
  );
  fifoFabOut_0 fifoFabOut_5(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_5 ),
       .io_deqData( fifoFabOut_5_io_deqData ),
       .io_enqRdy( fifoFabOut_5_io_enqRdy ),
       .io_deqRdy( T122 ),
       .io_enqValid( io_fabOutLocValid_5 ),
       .io_deqValid( fifoFabOut_5_io_deqValid ),
       .io_emptySpace( fifoFabOut_5_io_emptySpace ),
       .io_rst( T121 )
  );
  fifoFabOut_0 fifoFabOut_6(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_6 ),
       .io_deqData( fifoFabOut_6_io_deqData ),
       .io_enqRdy( fifoFabOut_6_io_enqRdy ),
       .io_deqRdy( T120 ),
       .io_enqValid( io_fabOutLocValid_6 ),
       .io_deqValid( fifoFabOut_6_io_deqValid ),
       .io_emptySpace( fifoFabOut_6_io_emptySpace ),
       .io_rst( T119 )
  );
  fifoFabOut_0 fifoFabOut_7(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_7 ),
       .io_deqData( fifoFabOut_7_io_deqData ),
       .io_enqRdy( fifoFabOut_7_io_enqRdy ),
       .io_deqRdy( T118 ),
       .io_enqValid( io_fabOutLocValid_7 ),
       .io_deqValid( fifoFabOut_7_io_deqValid ),
       .io_emptySpace( fifoFabOut_7_io_emptySpace ),
       .io_rst( T117 )
  );
  fifoFabOut_0 fifoFabOut_8(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_8 ),
       .io_deqData( fifoFabOut_8_io_deqData ),
       .io_enqRdy( fifoFabOut_8_io_enqRdy ),
       .io_deqRdy( T116 ),
       .io_enqValid( io_fabOutLocValid_8 ),
       .io_deqValid( fifoFabOut_8_io_deqValid ),
       .io_emptySpace( fifoFabOut_8_io_emptySpace ),
       .io_rst( T115 )
  );
  fifoFabOut_0 fifoFabOut_9(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_9 ),
       .io_deqData( fifoFabOut_9_io_deqData ),
       .io_enqRdy( fifoFabOut_9_io_enqRdy ),
       .io_deqRdy( T114 ),
       .io_enqValid( io_fabOutLocValid_9 ),
       .io_deqValid( fifoFabOut_9_io_deqValid ),
       .io_emptySpace( fifoFabOut_9_io_emptySpace ),
       .io_rst( T113 )
  );
  fifoFabOut_0 fifoFabOut_10(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_10 ),
       .io_deqData( fifoFabOut_10_io_deqData ),
       .io_enqRdy( fifoFabOut_10_io_enqRdy ),
       .io_deqRdy( T112 ),
       .io_enqValid( io_fabOutLocValid_10 ),
       .io_deqValid( fifoFabOut_10_io_deqValid ),
       .io_emptySpace( fifoFabOut_10_io_emptySpace ),
       .io_rst( T111 )
  );
  fifoFabOut_0 fifoFabOut_11(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_11 ),
       .io_deqData( fifoFabOut_11_io_deqData ),
       .io_enqRdy( fifoFabOut_11_io_enqRdy ),
       .io_deqRdy( T110 ),
       .io_enqValid( io_fabOutLocValid_11 ),
       .io_deqValid( fifoFabOut_11_io_deqValid ),
       .io_emptySpace( fifoFabOut_11_io_emptySpace ),
       .io_rst( T109 )
  );
  fifoFabOut_0 fifoFabOut_12(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_12 ),
       .io_deqData( fifoFabOut_12_io_deqData ),
       .io_enqRdy( fifoFabOut_12_io_enqRdy ),
       .io_deqRdy( T108 ),
       .io_enqValid( io_fabOutLocValid_12 ),
       .io_deqValid( fifoFabOut_12_io_deqValid ),
       .io_emptySpace( fifoFabOut_12_io_emptySpace ),
       .io_rst( T107 )
  );
  fifoFabOut_0 fifoFabOut_13(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_13 ),
       .io_deqData( fifoFabOut_13_io_deqData ),
       .io_enqRdy( fifoFabOut_13_io_enqRdy ),
       .io_deqRdy( T106 ),
       .io_enqValid( io_fabOutLocValid_13 ),
       .io_deqValid( fifoFabOut_13_io_deqValid ),
       .io_emptySpace( fifoFabOut_13_io_emptySpace ),
       .io_rst( T105 )
  );
  fifoFabOut_0 fifoFabOut_14(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_14 ),
       .io_deqData( fifoFabOut_14_io_deqData ),
       .io_enqRdy( fifoFabOut_14_io_enqRdy ),
       .io_deqRdy( T104 ),
       .io_enqValid( io_fabOutLocValid_14 ),
       .io_deqValid( fifoFabOut_14_io_deqValid ),
       .io_emptySpace( fifoFabOut_14_io_emptySpace ),
       .io_rst( T103 )
  );
  fifoFabOut_0 fifoFabOut_15(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_15 ),
       .io_deqData( fifoFabOut_15_io_deqData ),
       .io_enqRdy( fifoFabOut_15_io_enqRdy ),
       .io_deqRdy( T102 ),
       .io_enqValid( io_fabOutLocValid_15 ),
       .io_deqValid( fifoFabOut_15_io_deqValid ),
       .io_emptySpace( fifoFabOut_15_io_emptySpace ),
       .io_rst( T101 )
  );
  fifoFabOut_0 fifoFabOut_16(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_16 ),
       .io_deqData( fifoFabOut_16_io_deqData ),
       .io_enqRdy( fifoFabOut_16_io_enqRdy ),
       .io_deqRdy( T100 ),
       .io_enqValid( io_fabOutLocValid_16 ),
       .io_deqValid( fifoFabOut_16_io_deqValid ),
       .io_emptySpace( fifoFabOut_16_io_emptySpace ),
       .io_rst( T99 )
  );
  fifoFabOut_0 fifoFabOut_17(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_17 ),
       .io_deqData( fifoFabOut_17_io_deqData ),
       .io_enqRdy( fifoFabOut_17_io_enqRdy ),
       .io_deqRdy( T98 ),
       .io_enqValid( io_fabOutLocValid_17 ),
       .io_deqValid( fifoFabOut_17_io_deqValid ),
       .io_emptySpace( fifoFabOut_17_io_emptySpace ),
       .io_rst( T97 )
  );
  fifoFabOut_0 fifoFabOut_18(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_18 ),
       .io_deqData( fifoFabOut_18_io_deqData ),
       .io_enqRdy( fifoFabOut_18_io_enqRdy ),
       .io_deqRdy( T96 ),
       .io_enqValid( io_fabOutLocValid_18 ),
       .io_deqValid( fifoFabOut_18_io_deqValid ),
       .io_emptySpace( fifoFabOut_18_io_emptySpace ),
       .io_rst( T95 )
  );
  fifoFabOut_0 fifoFabOut_19(.clk(clk), .reset(reset),
       .io_enqData( io_fabOutLoc_19 ),
       .io_deqData( fifoFabOut_19_io_deqData ),
       .io_enqRdy( fifoFabOut_19_io_enqRdy ),
       .io_deqRdy( T94 ),
       .io_enqValid( io_fabOutLocValid_19 ),
       .io_deqValid( fifoFabOut_19_io_deqValid ),
       .io_emptySpace( fifoFabOut_19_io_emptySpace ),
       .io_rst( T93 )
  );
  fifoFabOut_1 outFifo(.clk(clk), .reset(reset),
       .io_enqData( T64 ),
       .io_deqData( outFifo_io_deqData ),
       .io_enqRdy( outFifo_io_enqRdy ),
       .io_deqRdy( io_locStoreRdy ),
       .io_enqValid( T1 ),
       .io_deqValid( outFifo_io_deqValid ),
       .io_emptySpace( outFifo_io_emptySpace ),
       .io_rst( T0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      muxValidReg_0 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_0 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_0 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_0 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_0 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_0 <= 1'h0;
    end else if(grantReg_3) begin
      muxValidReg_0 <= fifoFabOut_3_io_deqValid;
    end else if(grantReg_2) begin
      muxValidReg_0 <= fifoFabOut_2_io_deqValid;
    end else if(grantReg_1) begin
      muxValidReg_0 <= fifoFabOut_1_io_deqValid;
    end else if(grantReg_0) begin
      muxValidReg_0 <= fifoFabOut_io_deqValid;
    end
    if(reset) begin
      grantReg_0 <= 1'h0;
    end else begin
      grantReg_0 <= grantWire_0;
    end
    if(reset) begin
      grantReg_1 <= 1'h0;
    end else begin
      grantReg_1 <= grantWire_1;
    end
    if(reset) begin
      grantReg_2 <= 1'h0;
    end else begin
      grantReg_2 <= grantWire_2;
    end
    if(reset) begin
      grantReg_3 <= 1'h0;
    end else begin
      grantReg_3 <= grantWire_3;
    end
    if(reset) begin
      muxValidReg_1 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_1 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_1 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_1 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_1 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_1 <= 1'h0;
    end else if(grantReg_7) begin
      muxValidReg_1 <= fifoFabOut_7_io_deqValid;
    end else if(grantReg_6) begin
      muxValidReg_1 <= fifoFabOut_6_io_deqValid;
    end else if(grantReg_5) begin
      muxValidReg_1 <= fifoFabOut_5_io_deqValid;
    end else if(grantReg_4) begin
      muxValidReg_1 <= fifoFabOut_4_io_deqValid;
    end
    if(reset) begin
      grantReg_4 <= 1'h0;
    end else begin
      grantReg_4 <= grantWire_4;
    end
    if(reset) begin
      grantReg_5 <= 1'h0;
    end else begin
      grantReg_5 <= grantWire_5;
    end
    if(reset) begin
      grantReg_6 <= 1'h0;
    end else begin
      grantReg_6 <= grantWire_6;
    end
    if(reset) begin
      grantReg_7 <= 1'h0;
    end else begin
      grantReg_7 <= grantWire_7;
    end
    if(reset) begin
      muxValidReg_2 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_2 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_2 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_2 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_2 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_2 <= 1'h0;
    end else if(grantReg_11) begin
      muxValidReg_2 <= fifoFabOut_11_io_deqValid;
    end else if(grantReg_10) begin
      muxValidReg_2 <= fifoFabOut_10_io_deqValid;
    end else if(grantReg_9) begin
      muxValidReg_2 <= fifoFabOut_9_io_deqValid;
    end else if(grantReg_8) begin
      muxValidReg_2 <= fifoFabOut_8_io_deqValid;
    end
    if(reset) begin
      grantReg_8 <= 1'h0;
    end else begin
      grantReg_8 <= grantWire_8;
    end
    if(reset) begin
      grantReg_9 <= 1'h0;
    end else begin
      grantReg_9 <= grantWire_9;
    end
    if(reset) begin
      grantReg_10 <= 1'h0;
    end else begin
      grantReg_10 <= grantWire_10;
    end
    if(reset) begin
      grantReg_11 <= 1'h0;
    end else begin
      grantReg_11 <= grantWire_11;
    end
    if(reset) begin
      muxValidReg_3 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_3 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_3 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_3 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_3 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_3 <= 1'h0;
    end else if(grantReg_15) begin
      muxValidReg_3 <= fifoFabOut_15_io_deqValid;
    end else if(grantReg_14) begin
      muxValidReg_3 <= fifoFabOut_14_io_deqValid;
    end else if(grantReg_13) begin
      muxValidReg_3 <= fifoFabOut_13_io_deqValid;
    end else if(grantReg_12) begin
      muxValidReg_3 <= fifoFabOut_12_io_deqValid;
    end
    if(reset) begin
      grantReg_12 <= 1'h0;
    end else begin
      grantReg_12 <= grantWire_12;
    end
    if(reset) begin
      grantReg_13 <= 1'h0;
    end else begin
      grantReg_13 <= grantWire_13;
    end
    if(reset) begin
      grantReg_14 <= 1'h0;
    end else begin
      grantReg_14 <= grantWire_14;
    end
    if(reset) begin
      grantReg_15 <= 1'h0;
    end else begin
      grantReg_15 <= grantWire_15;
    end
    if(reset) begin
      muxValidReg_4 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_4 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_4 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_4 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_4 <= 1'h0;
    end else if(io_rst) begin
      muxValidReg_4 <= 1'h0;
    end else if(grantReg_19) begin
      muxValidReg_4 <= fifoFabOut_19_io_deqValid;
    end else if(grantReg_18) begin
      muxValidReg_4 <= fifoFabOut_18_io_deqValid;
    end else if(grantReg_17) begin
      muxValidReg_4 <= fifoFabOut_17_io_deqValid;
    end else if(grantReg_16) begin
      muxValidReg_4 <= fifoFabOut_16_io_deqValid;
    end
    if(reset) begin
      grantReg_16 <= 1'h0;
    end else begin
      grantReg_16 <= grantWire_16;
    end
    if(reset) begin
      grantReg_17 <= 1'h0;
    end else begin
      grantReg_17 <= grantWire_17;
    end
    if(reset) begin
      grantReg_18 <= 1'h0;
    end else begin
      grantReg_18 <= grantWire_18;
    end
    if(reset) begin
      grantReg_19 <= 1'h0;
    end else begin
      grantReg_19 <= grantWire_19;
    end
    if(reset) begin
      muxReg_0 <= 56'h0;
    end else if(grantReg_3) begin
      muxReg_0 <= fifoFabOut_3_io_deqData;
    end else if(grantReg_2) begin
      muxReg_0 <= fifoFabOut_2_io_deqData;
    end else if(grantReg_1) begin
      muxReg_0 <= fifoFabOut_1_io_deqData;
    end else if(grantReg_0) begin
      muxReg_0 <= fifoFabOut_io_deqData;
    end
    if(reset) begin
      muxReg_1 <= 56'h0;
    end else if(grantReg_7) begin
      muxReg_1 <= fifoFabOut_7_io_deqData;
    end else if(grantReg_6) begin
      muxReg_1 <= fifoFabOut_6_io_deqData;
    end else if(grantReg_5) begin
      muxReg_1 <= fifoFabOut_5_io_deqData;
    end else if(grantReg_4) begin
      muxReg_1 <= fifoFabOut_4_io_deqData;
    end
    if(reset) begin
      muxReg_2 <= 56'h0;
    end else if(grantReg_11) begin
      muxReg_2 <= fifoFabOut_11_io_deqData;
    end else if(grantReg_10) begin
      muxReg_2 <= fifoFabOut_10_io_deqData;
    end else if(grantReg_9) begin
      muxReg_2 <= fifoFabOut_9_io_deqData;
    end else if(grantReg_8) begin
      muxReg_2 <= fifoFabOut_8_io_deqData;
    end
    if(reset) begin
      muxReg_3 <= 56'h0;
    end else if(grantReg_15) begin
      muxReg_3 <= fifoFabOut_15_io_deqData;
    end else if(grantReg_14) begin
      muxReg_3 <= fifoFabOut_14_io_deqData;
    end else if(grantReg_13) begin
      muxReg_3 <= fifoFabOut_13_io_deqData;
    end else if(grantReg_12) begin
      muxReg_3 <= fifoFabOut_12_io_deqData;
    end
    if(reset) begin
      muxReg_4 <= 56'h0;
    end else if(grantReg_19) begin
      muxReg_4 <= fifoFabOut_19_io_deqData;
    end else if(grantReg_18) begin
      muxReg_4 <= fifoFabOut_18_io_deqData;
    end else if(grantReg_17) begin
      muxReg_4 <= fifoFabOut_17_io_deqData;
    end else if(grantReg_16) begin
      muxReg_4 <= fifoFabOut_16_io_deqData;
    end
  end
endmodule

module fabOutSeqTop(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input [31:0] io_fabOut_19,
    input [31:0] io_fabOut_18,
    input [31:0] io_fabOut_17,
    input [31:0] io_fabOut_16,
    input [31:0] io_fabOut_15,
    input [31:0] io_fabOut_14,
    input [31:0] io_fabOut_13,
    input [31:0] io_fabOut_12,
    input [31:0] io_fabOut_11,
    input [31:0] io_fabOut_10,
    input [31:0] io_fabOut_9,
    input [31:0] io_fabOut_8,
    input [31:0] io_fabOut_7,
    input [31:0] io_fabOut_6,
    input [31:0] io_fabOut_5,
    input [31:0] io_fabOut_4,
    input [31:0] io_fabOut_3,
    input [31:0] io_fabOut_2,
    input [31:0] io_fabOut_1,
    input [31:0] io_fabOut_0,
    input  io_fabOutValid_19,
    input  io_fabOutValid_18,
    input  io_fabOutValid_17,
    input  io_fabOutValid_16,
    input  io_fabOutValid_15,
    input  io_fabOutValid_14,
    input  io_fabOutValid_13,
    input  io_fabOutValid_12,
    input  io_fabOutValid_11,
    input  io_fabOutValid_10,
    input  io_fabOutValid_9,
    input  io_fabOutValid_8,
    input  io_fabOutValid_7,
    input  io_fabOutValid_6,
    input  io_fabOutValid_5,
    input  io_fabOutValid_4,
    input  io_fabOutValid_3,
    input  io_fabOutValid_2,
    input  io_fabOutValid_1,
    input  io_fabOutValid_0,
    output io_fabOutRdy_19,
    output io_fabOutRdy_18,
    output io_fabOutRdy_17,
    output io_fabOutRdy_16,
    output io_fabOutRdy_15,
    output io_fabOutRdy_14,
    output io_fabOutRdy_13,
    output io_fabOutRdy_12,
    output io_fabOutRdy_11,
    output io_fabOutRdy_10,
    output io_fabOutRdy_9,
    output io_fabOutRdy_8,
    output io_fabOutRdy_7,
    output io_fabOutRdy_6,
    output io_fabOutRdy_5,
    output io_fabOutRdy_4,
    output io_fabOutRdy_3,
    output io_fabOutRdy_2,
    output io_fabOutRdy_1,
    output io_fabOutRdy_0,
    output[31:0] io_fabOutStore_19,
    output[31:0] io_fabOutStore_18,
    output[31:0] io_fabOutStore_17,
    output[31:0] io_fabOutStore_16,
    output[31:0] io_fabOutStore_15,
    output[31:0] io_fabOutStore_14,
    output[31:0] io_fabOutStore_13,
    output[31:0] io_fabOutStore_12,
    output[31:0] io_fabOutStore_11,
    output[31:0] io_fabOutStore_10,
    output[31:0] io_fabOutStore_9,
    output[31:0] io_fabOutStore_8,
    output[31:0] io_fabOutStore_7,
    output[31:0] io_fabOutStore_6,
    output[31:0] io_fabOutStore_5,
    output[31:0] io_fabOutStore_4,
    output[31:0] io_fabOutStore_3,
    output[31:0] io_fabOutStore_2,
    output[31:0] io_fabOutStore_1,
    output[31:0] io_fabOutStore_0,
    output io_fabOutStoreValid_19,
    output io_fabOutStoreValid_18,
    output io_fabOutStoreValid_17,
    output io_fabOutStoreValid_16,
    output io_fabOutStoreValid_15,
    output io_fabOutStoreValid_14,
    output io_fabOutStoreValid_13,
    output io_fabOutStoreValid_12,
    output io_fabOutStoreValid_11,
    output io_fabOutStoreValid_10,
    output io_fabOutStoreValid_9,
    output io_fabOutStoreValid_8,
    output io_fabOutStoreValid_7,
    output io_fabOutStoreValid_6,
    output io_fabOutStoreValid_5,
    output io_fabOutStoreValid_4,
    output io_fabOutStoreValid_3,
    output io_fabOutStoreValid_2,
    output io_fabOutStoreValid_1,
    output io_fabOutStoreValid_0,
    input  io_fabOutStoreRdy_19,
    input  io_fabOutStoreRdy_18,
    input  io_fabOutStoreRdy_17,
    input  io_fabOutStoreRdy_16,
    input  io_fabOutStoreRdy_15,
    input  io_fabOutStoreRdy_14,
    input  io_fabOutStoreRdy_13,
    input  io_fabOutStoreRdy_12,
    input  io_fabOutStoreRdy_11,
    input  io_fabOutStoreRdy_10,
    input  io_fabOutStoreRdy_9,
    input  io_fabOutStoreRdy_8,
    input  io_fabOutStoreRdy_7,
    input  io_fabOutStoreRdy_6,
    input  io_fabOutStoreRdy_5,
    input  io_fabOutStoreRdy_4,
    input  io_fabOutStoreRdy_3,
    input  io_fabOutStoreRdy_2,
    input  io_fabOutStoreRdy_1,
    input  io_fabOutStoreRdy_0,
    output[87:0] io_fabOutLoc_7,
    output[87:0] io_fabOutLoc_6,
    output[87:0] io_fabOutLoc_5,
    output[87:0] io_fabOutLoc_4,
    output[87:0] io_fabOutLoc_3,
    output[87:0] io_fabOutLoc_2,
    output[87:0] io_fabOutLoc_1,
    output[87:0] io_fabOutLoc_0,
    output io_fabOutLocValid_7,
    output io_fabOutLocValid_6,
    output io_fabOutLocValid_5,
    output io_fabOutLocValid_4,
    output io_fabOutLocValid_3,
    output io_fabOutLocValid_2,
    output io_fabOutLocValid_1,
    output io_fabOutLocValid_0,
    input  io_fabOutLocRdy_7,
    input  io_fabOutLocRdy_6,
    input  io_fabOutLocRdy_5,
    input  io_fabOutLocRdy_4,
    input  io_fabOutLocRdy_3,
    input  io_fabOutLocRdy_2,
    input  io_fabOutLocRdy_1,
    input  io_fabOutLocRdy_0
);

  wire[55:0] T0;
  wire[55:0] T1;
  wire[55:0] T2;
  wire[55:0] T3;
  wire[55:0] T4;
  wire[55:0] T5;
  wire[55:0] T6;
  wire[55:0] T7;
  wire[55:0] T8;
  wire[55:0] T9;
  wire[55:0] T10;
  wire[55:0] T11;
  wire[55:0] T12;
  wire[55:0] T13;
  wire[55:0] T14;
  wire[55:0] T15;
  wire[55:0] T16;
  wire[55:0] T17;
  wire[55:0] T18;
  wire[55:0] T19;
  wire[55:0] T20;
  wire[55:0] T21;
  wire[55:0] T22;
  wire[55:0] T23;
  wire[55:0] T24;
  wire[55:0] T25;
  wire[55:0] T26;
  wire[55:0] T27;
  wire[55:0] T28;
  wire[55:0] T29;
  wire[55:0] T30;
  wire[55:0] T31;
  wire[55:0] T32;
  wire[55:0] T33;
  wire[55:0] T34;
  wire[55:0] T35;
  wire[55:0] T36;
  wire[55:0] T37;
  wire[55:0] T38;
  wire[55:0] T39;
  wire[55:0] T40;
  wire[55:0] T41;
  wire[55:0] T42;
  wire[55:0] T43;
  wire[55:0] T44;
  wire[55:0] T45;
  wire[55:0] T46;
  wire[55:0] T47;
  wire[55:0] T48;
  wire[55:0] T49;
  wire[55:0] T50;
  wire[55:0] T51;
  wire[55:0] T52;
  wire[55:0] T53;
  wire[55:0] T54;
  wire[55:0] T55;
  wire[55:0] T56;
  wire[55:0] T57;
  wire[55:0] T58;
  wire[55:0] T59;
  wire[55:0] T60;
  wire[55:0] T61;
  wire[55:0] T62;
  wire[55:0] T63;
  wire[55:0] T64;
  wire[55:0] T65;
  wire[55:0] T66;
  wire[55:0] T67;
  wire[55:0] T68;
  wire[55:0] T69;
  wire[55:0] T70;
  wire[55:0] T71;
  wire[55:0] T72;
  wire[55:0] T73;
  wire[55:0] T74;
  wire[55:0] T75;
  wire[55:0] T76;
  wire[55:0] T77;
  wire[55:0] T78;
  wire[55:0] T79;
  wire[55:0] T80;
  wire[55:0] T81;
  wire[55:0] T82;
  wire[55:0] T83;
  wire[55:0] T84;
  wire[55:0] T85;
  wire[55:0] T86;
  wire[55:0] T87;
  wire[55:0] T88;
  wire[55:0] T89;
  wire[55:0] T90;
  wire[55:0] T91;
  wire[55:0] T92;
  wire[55:0] T93;
  wire[55:0] T94;
  wire[55:0] T95;
  wire[55:0] T96;
  wire[55:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[55:0] T100;
  wire[55:0] T101;
  wire[55:0] T102;
  wire[55:0] T103;
  wire[55:0] T104;
  wire[55:0] T105;
  wire[55:0] T106;
  wire[55:0] T107;
  wire[55:0] T108;
  wire[55:0] T109;
  wire[55:0] T110;
  wire[55:0] T111;
  wire[55:0] T112;
  wire[55:0] T113;
  wire[55:0] T114;
  wire[55:0] T115;
  wire[55:0] T116;
  wire[55:0] T117;
  wire[55:0] T118;
  wire[55:0] T119;
  wire[55:0] T120;
  wire[55:0] T121;
  wire[55:0] T122;
  wire[55:0] T123;
  wire[55:0] T124;
  wire[55:0] T125;
  wire[55:0] T126;
  wire[55:0] T127;
  wire[55:0] T128;
  wire[55:0] T129;
  wire[55:0] T130;
  wire[55:0] T131;
  wire[55:0] T132;
  wire[55:0] T133;
  wire[55:0] T134;
  wire[55:0] T135;
  wire[55:0] T136;
  wire[55:0] T137;
  wire[55:0] T138;
  wire[55:0] T139;
  wire[55:0] T140;
  wire[55:0] T141;
  wire[55:0] T142;
  wire[55:0] T143;
  wire[55:0] T144;
  wire[55:0] T145;
  wire[55:0] T146;
  wire[55:0] T147;
  wire[55:0] T148;
  wire[55:0] T149;
  wire[55:0] T150;
  wire[55:0] T151;
  wire[55:0] T152;
  wire[55:0] T153;
  wire[55:0] T154;
  wire[55:0] T155;
  wire[55:0] T156;
  wire[55:0] T157;
  wire[55:0] T158;
  wire[55:0] T159;
  wire[87:0] T160;
  wire[87:0] T161;
  wire[87:0] T162;
  wire[87:0] T163;
  wire[87:0] T164;
  wire[87:0] T165;
  wire[87:0] T166;
  wire[87:0] T167;
  wire[55:0] fabOutSeqArb_io_locStoreData;
  wire fabOutSeqArb_io_locStoreValid;
  wire[55:0] fabOutSeqArb_1_io_locStoreData;
  wire fabOutSeqArb_1_io_locStoreValid;
  wire[55:0] fabOutSeqArb_2_io_locStoreData;
  wire fabOutSeqArb_2_io_locStoreValid;
  wire[55:0] fabOutSeqArb_3_io_locStoreData;
  wire fabOutSeqArb_3_io_locStoreValid;
  wire[55:0] fabOutSeqArb_4_io_locStoreData;
  wire fabOutSeqArb_4_io_locStoreValid;
  wire[55:0] fabOutSeqArb_5_io_locStoreData;
  wire fabOutSeqArb_5_io_locStoreValid;
  wire[55:0] fabOutSeqArb_6_io_locStoreData;
  wire fabOutSeqArb_6_io_locStoreValid;
  wire fabOutSeqArb_7_io_fabOutLocRdy_19;
  wire fabOutSeqArb_7_io_fabOutLocRdy_18;
  wire fabOutSeqArb_7_io_fabOutLocRdy_17;
  wire fabOutSeqArb_7_io_fabOutLocRdy_16;
  wire fabOutSeqArb_7_io_fabOutLocRdy_15;
  wire fabOutSeqArb_7_io_fabOutLocRdy_14;
  wire fabOutSeqArb_7_io_fabOutLocRdy_13;
  wire fabOutSeqArb_7_io_fabOutLocRdy_12;
  wire fabOutSeqArb_7_io_fabOutLocRdy_11;
  wire fabOutSeqArb_7_io_fabOutLocRdy_10;
  wire fabOutSeqArb_7_io_fabOutLocRdy_9;
  wire fabOutSeqArb_7_io_fabOutLocRdy_8;
  wire fabOutSeqArb_7_io_fabOutLocRdy_7;
  wire fabOutSeqArb_7_io_fabOutLocRdy_6;
  wire fabOutSeqArb_7_io_fabOutLocRdy_5;
  wire fabOutSeqArb_7_io_fabOutLocRdy_4;
  wire fabOutSeqArb_7_io_fabOutLocRdy_3;
  wire fabOutSeqArb_7_io_fabOutLocRdy_2;
  wire fabOutSeqArb_7_io_fabOutLocRdy_1;
  wire fabOutSeqArb_7_io_fabOutLocRdy_0;
  wire[55:0] fabOutSeqArb_7_io_locStoreData;
  wire fabOutSeqArb_7_io_locStoreValid;
  wire fabOutSeqIntClass_io_fabOutRdy_19;
  wire fabOutSeqIntClass_io_fabOutRdy_18;
  wire fabOutSeqIntClass_io_fabOutRdy_17;
  wire fabOutSeqIntClass_io_fabOutRdy_16;
  wire fabOutSeqIntClass_io_fabOutRdy_15;
  wire fabOutSeqIntClass_io_fabOutRdy_14;
  wire fabOutSeqIntClass_io_fabOutRdy_13;
  wire fabOutSeqIntClass_io_fabOutRdy_12;
  wire fabOutSeqIntClass_io_fabOutRdy_11;
  wire fabOutSeqIntClass_io_fabOutRdy_10;
  wire fabOutSeqIntClass_io_fabOutRdy_9;
  wire fabOutSeqIntClass_io_fabOutRdy_8;
  wire fabOutSeqIntClass_io_fabOutRdy_7;
  wire fabOutSeqIntClass_io_fabOutRdy_6;
  wire fabOutSeqIntClass_io_fabOutRdy_5;
  wire fabOutSeqIntClass_io_fabOutRdy_4;
  wire fabOutSeqIntClass_io_fabOutRdy_3;
  wire fabOutSeqIntClass_io_fabOutRdy_2;
  wire fabOutSeqIntClass_io_fabOutRdy_1;
  wire fabOutSeqIntClass_io_fabOutRdy_0;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_19;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_18;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_17;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_16;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_15;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_14;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_13;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_12;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_11;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_10;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_9;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_8;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_7;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_6;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_5;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_4;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_3;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_2;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_1;
  wire[31:0] fabOutSeqIntClass_io_fabOutStore_0;
  wire fabOutSeqIntClass_io_fabOutStoreValid_19;
  wire fabOutSeqIntClass_io_fabOutStoreValid_18;
  wire fabOutSeqIntClass_io_fabOutStoreValid_17;
  wire fabOutSeqIntClass_io_fabOutStoreValid_16;
  wire fabOutSeqIntClass_io_fabOutStoreValid_15;
  wire fabOutSeqIntClass_io_fabOutStoreValid_14;
  wire fabOutSeqIntClass_io_fabOutStoreValid_13;
  wire fabOutSeqIntClass_io_fabOutStoreValid_12;
  wire fabOutSeqIntClass_io_fabOutStoreValid_11;
  wire fabOutSeqIntClass_io_fabOutStoreValid_10;
  wire fabOutSeqIntClass_io_fabOutStoreValid_9;
  wire fabOutSeqIntClass_io_fabOutStoreValid_8;
  wire fabOutSeqIntClass_io_fabOutStoreValid_7;
  wire fabOutSeqIntClass_io_fabOutStoreValid_6;
  wire fabOutSeqIntClass_io_fabOutStoreValid_5;
  wire fabOutSeqIntClass_io_fabOutStoreValid_4;
  wire fabOutSeqIntClass_io_fabOutStoreValid_3;
  wire fabOutSeqIntClass_io_fabOutStoreValid_2;
  wire fabOutSeqIntClass_io_fabOutStoreValid_1;
  wire fabOutSeqIntClass_io_fabOutStoreValid_0;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_19;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_18;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_17;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_16;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_15;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_14;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_13;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_12;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_11;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_10;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_9;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_8;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_7;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_6;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_5;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_4;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_3;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_2;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_1;
  wire[87:0] fabOutSeqIntClass_io_fabOutLoc_0;
  wire fabOutSeqIntClass_io_fabOutLocValid_19;
  wire fabOutSeqIntClass_io_fabOutLocValid_18;
  wire fabOutSeqIntClass_io_fabOutLocValid_17;
  wire fabOutSeqIntClass_io_fabOutLocValid_16;
  wire fabOutSeqIntClass_io_fabOutLocValid_15;
  wire fabOutSeqIntClass_io_fabOutLocValid_14;
  wire fabOutSeqIntClass_io_fabOutLocValid_13;
  wire fabOutSeqIntClass_io_fabOutLocValid_12;
  wire fabOutSeqIntClass_io_fabOutLocValid_11;
  wire fabOutSeqIntClass_io_fabOutLocValid_10;
  wire fabOutSeqIntClass_io_fabOutLocValid_9;
  wire fabOutSeqIntClass_io_fabOutLocValid_8;
  wire fabOutSeqIntClass_io_fabOutLocValid_7;
  wire fabOutSeqIntClass_io_fabOutLocValid_6;
  wire fabOutSeqIntClass_io_fabOutLocValid_5;
  wire fabOutSeqIntClass_io_fabOutLocValid_4;
  wire fabOutSeqIntClass_io_fabOutLocValid_3;
  wire fabOutSeqIntClass_io_fabOutLocValid_2;
  wire fabOutSeqIntClass_io_fabOutLocValid_1;
  wire fabOutSeqIntClass_io_fabOutLocValid_0;
  wire fabOutSeqIntClass_io_rst;


  assign T0 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T1 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T2 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T3 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T4 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T5 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T6 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T7 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T8 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T9 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T10 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T11 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T12 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T13 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T14 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T15 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T16 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T17 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T18 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T19 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T20 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T21 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T22 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T23 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T24 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T25 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T26 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T27 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T28 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T29 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T30 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T31 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T32 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T33 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T34 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T35 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T36 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T37 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T38 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T39 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T40 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T41 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T42 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T43 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T44 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T45 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T46 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T47 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T48 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T49 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T50 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T51 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T52 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T53 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T54 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T55 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T56 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T57 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T58 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T59 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T60 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T61 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T62 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T63 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T64 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T65 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T66 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T67 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T68 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T69 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T70 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T71 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T72 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T73 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T74 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T75 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T76 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T77 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T78 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T79 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T80 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T81 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T82 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T83 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T84 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T85 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T86 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T87 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T88 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T89 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T90 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T91 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T92 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T93 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T94 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T95 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T96 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T97 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T98 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T99 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T100 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T101 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T102 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T103 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T104 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T105 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T106 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T107 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T108 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T109 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T110 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T111 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T112 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T113 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T114 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T115 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T116 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T117 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T118 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T119 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T120 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T121 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T122 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T123 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T124 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T125 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T126 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T127 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T128 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T129 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T130 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T131 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T132 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T133 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T134 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T135 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T136 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T137 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T138 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T139 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign T140 = fabOutSeqIntClass_io_fabOutLoc_0[6'h37:1'h0];
  assign T141 = fabOutSeqIntClass_io_fabOutLoc_1[6'h37:1'h0];
  assign T142 = fabOutSeqIntClass_io_fabOutLoc_2[6'h37:1'h0];
  assign T143 = fabOutSeqIntClass_io_fabOutLoc_3[6'h37:1'h0];
  assign T144 = fabOutSeqIntClass_io_fabOutLoc_4[6'h37:1'h0];
  assign T145 = fabOutSeqIntClass_io_fabOutLoc_5[6'h37:1'h0];
  assign T146 = fabOutSeqIntClass_io_fabOutLoc_6[6'h37:1'h0];
  assign T147 = fabOutSeqIntClass_io_fabOutLoc_7[6'h37:1'h0];
  assign T148 = fabOutSeqIntClass_io_fabOutLoc_8[6'h37:1'h0];
  assign T149 = fabOutSeqIntClass_io_fabOutLoc_9[6'h37:1'h0];
  assign T150 = fabOutSeqIntClass_io_fabOutLoc_10[6'h37:1'h0];
  assign T151 = fabOutSeqIntClass_io_fabOutLoc_11[6'h37:1'h0];
  assign T152 = fabOutSeqIntClass_io_fabOutLoc_12[6'h37:1'h0];
  assign T153 = fabOutSeqIntClass_io_fabOutLoc_13[6'h37:1'h0];
  assign T154 = fabOutSeqIntClass_io_fabOutLoc_14[6'h37:1'h0];
  assign T155 = fabOutSeqIntClass_io_fabOutLoc_15[6'h37:1'h0];
  assign T156 = fabOutSeqIntClass_io_fabOutLoc_16[6'h37:1'h0];
  assign T157 = fabOutSeqIntClass_io_fabOutLoc_17[6'h37:1'h0];
  assign T158 = fabOutSeqIntClass_io_fabOutLoc_18[6'h37:1'h0];
  assign T159 = fabOutSeqIntClass_io_fabOutLoc_19[6'h37:1'h0];
  assign io_fabOutLocValid_0 = fabOutSeqArb_io_locStoreValid;
  assign io_fabOutLocValid_1 = fabOutSeqArb_1_io_locStoreValid;
  assign io_fabOutLocValid_2 = fabOutSeqArb_2_io_locStoreValid;
  assign io_fabOutLocValid_3 = fabOutSeqArb_3_io_locStoreValid;
  assign io_fabOutLocValid_4 = fabOutSeqArb_4_io_locStoreValid;
  assign io_fabOutLocValid_5 = fabOutSeqArb_5_io_locStoreValid;
  assign io_fabOutLocValid_6 = fabOutSeqArb_6_io_locStoreValid;
  assign io_fabOutLocValid_7 = fabOutSeqArb_7_io_locStoreValid;
  assign io_fabOutLoc_0 = T160;
  assign T160 = {32'h0, fabOutSeqArb_io_locStoreData};
  assign io_fabOutLoc_1 = T161;
  assign T161 = {32'h0, fabOutSeqArb_1_io_locStoreData};
  assign io_fabOutLoc_2 = T162;
  assign T162 = {32'h0, fabOutSeqArb_2_io_locStoreData};
  assign io_fabOutLoc_3 = T163;
  assign T163 = {32'h0, fabOutSeqArb_3_io_locStoreData};
  assign io_fabOutLoc_4 = T164;
  assign T164 = {32'h0, fabOutSeqArb_4_io_locStoreData};
  assign io_fabOutLoc_5 = T165;
  assign T165 = {32'h0, fabOutSeqArb_5_io_locStoreData};
  assign io_fabOutLoc_6 = T166;
  assign T166 = {32'h0, fabOutSeqArb_6_io_locStoreData};
  assign io_fabOutLoc_7 = T167;
  assign T167 = {32'h0, fabOutSeqArb_7_io_locStoreData};
  assign io_fabOutStoreValid_0 = fabOutSeqIntClass_io_fabOutStoreValid_0;
  assign io_fabOutStoreValid_1 = fabOutSeqIntClass_io_fabOutStoreValid_1;
  assign io_fabOutStoreValid_2 = fabOutSeqIntClass_io_fabOutStoreValid_2;
  assign io_fabOutStoreValid_3 = fabOutSeqIntClass_io_fabOutStoreValid_3;
  assign io_fabOutStoreValid_4 = fabOutSeqIntClass_io_fabOutStoreValid_4;
  assign io_fabOutStoreValid_5 = fabOutSeqIntClass_io_fabOutStoreValid_5;
  assign io_fabOutStoreValid_6 = fabOutSeqIntClass_io_fabOutStoreValid_6;
  assign io_fabOutStoreValid_7 = fabOutSeqIntClass_io_fabOutStoreValid_7;
  assign io_fabOutStoreValid_8 = fabOutSeqIntClass_io_fabOutStoreValid_8;
  assign io_fabOutStoreValid_9 = fabOutSeqIntClass_io_fabOutStoreValid_9;
  assign io_fabOutStoreValid_10 = fabOutSeqIntClass_io_fabOutStoreValid_10;
  assign io_fabOutStoreValid_11 = fabOutSeqIntClass_io_fabOutStoreValid_11;
  assign io_fabOutStoreValid_12 = fabOutSeqIntClass_io_fabOutStoreValid_12;
  assign io_fabOutStoreValid_13 = fabOutSeqIntClass_io_fabOutStoreValid_13;
  assign io_fabOutStoreValid_14 = fabOutSeqIntClass_io_fabOutStoreValid_14;
  assign io_fabOutStoreValid_15 = fabOutSeqIntClass_io_fabOutStoreValid_15;
  assign io_fabOutStoreValid_16 = fabOutSeqIntClass_io_fabOutStoreValid_16;
  assign io_fabOutStoreValid_17 = fabOutSeqIntClass_io_fabOutStoreValid_17;
  assign io_fabOutStoreValid_18 = fabOutSeqIntClass_io_fabOutStoreValid_18;
  assign io_fabOutStoreValid_19 = fabOutSeqIntClass_io_fabOutStoreValid_19;
  assign io_fabOutStore_0 = fabOutSeqIntClass_io_fabOutStore_0;
  assign io_fabOutStore_1 = fabOutSeqIntClass_io_fabOutStore_1;
  assign io_fabOutStore_2 = fabOutSeqIntClass_io_fabOutStore_2;
  assign io_fabOutStore_3 = fabOutSeqIntClass_io_fabOutStore_3;
  assign io_fabOutStore_4 = fabOutSeqIntClass_io_fabOutStore_4;
  assign io_fabOutStore_5 = fabOutSeqIntClass_io_fabOutStore_5;
  assign io_fabOutStore_6 = fabOutSeqIntClass_io_fabOutStore_6;
  assign io_fabOutStore_7 = fabOutSeqIntClass_io_fabOutStore_7;
  assign io_fabOutStore_8 = fabOutSeqIntClass_io_fabOutStore_8;
  assign io_fabOutStore_9 = fabOutSeqIntClass_io_fabOutStore_9;
  assign io_fabOutStore_10 = fabOutSeqIntClass_io_fabOutStore_10;
  assign io_fabOutStore_11 = fabOutSeqIntClass_io_fabOutStore_11;
  assign io_fabOutStore_12 = fabOutSeqIntClass_io_fabOutStore_12;
  assign io_fabOutStore_13 = fabOutSeqIntClass_io_fabOutStore_13;
  assign io_fabOutStore_14 = fabOutSeqIntClass_io_fabOutStore_14;
  assign io_fabOutStore_15 = fabOutSeqIntClass_io_fabOutStore_15;
  assign io_fabOutStore_16 = fabOutSeqIntClass_io_fabOutStore_16;
  assign io_fabOutStore_17 = fabOutSeqIntClass_io_fabOutStore_17;
  assign io_fabOutStore_18 = fabOutSeqIntClass_io_fabOutStore_18;
  assign io_fabOutStore_19 = fabOutSeqIntClass_io_fabOutStore_19;
  assign io_fabOutRdy_0 = fabOutSeqIntClass_io_fabOutRdy_0;
  assign io_fabOutRdy_1 = fabOutSeqIntClass_io_fabOutRdy_1;
  assign io_fabOutRdy_2 = fabOutSeqIntClass_io_fabOutRdy_2;
  assign io_fabOutRdy_3 = fabOutSeqIntClass_io_fabOutRdy_3;
  assign io_fabOutRdy_4 = fabOutSeqIntClass_io_fabOutRdy_4;
  assign io_fabOutRdy_5 = fabOutSeqIntClass_io_fabOutRdy_5;
  assign io_fabOutRdy_6 = fabOutSeqIntClass_io_fabOutRdy_6;
  assign io_fabOutRdy_7 = fabOutSeqIntClass_io_fabOutRdy_7;
  assign io_fabOutRdy_8 = fabOutSeqIntClass_io_fabOutRdy_8;
  assign io_fabOutRdy_9 = fabOutSeqIntClass_io_fabOutRdy_9;
  assign io_fabOutRdy_10 = fabOutSeqIntClass_io_fabOutRdy_10;
  assign io_fabOutRdy_11 = fabOutSeqIntClass_io_fabOutRdy_11;
  assign io_fabOutRdy_12 = fabOutSeqIntClass_io_fabOutRdy_12;
  assign io_fabOutRdy_13 = fabOutSeqIntClass_io_fabOutRdy_13;
  assign io_fabOutRdy_14 = fabOutSeqIntClass_io_fabOutRdy_14;
  assign io_fabOutRdy_15 = fabOutSeqIntClass_io_fabOutRdy_15;
  assign io_fabOutRdy_16 = fabOutSeqIntClass_io_fabOutRdy_16;
  assign io_fabOutRdy_17 = fabOutSeqIntClass_io_fabOutRdy_17;
  assign io_fabOutRdy_18 = fabOutSeqIntClass_io_fabOutRdy_18;
  assign io_fabOutRdy_19 = fabOutSeqIntClass_io_fabOutRdy_19;
  fabOutSeq fabOutSeqIntClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_fabOut_19( io_fabOut_19 ),
       .io_fabOut_18( io_fabOut_18 ),
       .io_fabOut_17( io_fabOut_17 ),
       .io_fabOut_16( io_fabOut_16 ),
       .io_fabOut_15( io_fabOut_15 ),
       .io_fabOut_14( io_fabOut_14 ),
       .io_fabOut_13( io_fabOut_13 ),
       .io_fabOut_12( io_fabOut_12 ),
       .io_fabOut_11( io_fabOut_11 ),
       .io_fabOut_10( io_fabOut_10 ),
       .io_fabOut_9( io_fabOut_9 ),
       .io_fabOut_8( io_fabOut_8 ),
       .io_fabOut_7( io_fabOut_7 ),
       .io_fabOut_6( io_fabOut_6 ),
       .io_fabOut_5( io_fabOut_5 ),
       .io_fabOut_4( io_fabOut_4 ),
       .io_fabOut_3( io_fabOut_3 ),
       .io_fabOut_2( io_fabOut_2 ),
       .io_fabOut_1( io_fabOut_1 ),
       .io_fabOut_0( io_fabOut_0 ),
       .io_fabOutValid_19( io_fabOutValid_19 ),
       .io_fabOutValid_18( io_fabOutValid_18 ),
       .io_fabOutValid_17( io_fabOutValid_17 ),
       .io_fabOutValid_16( io_fabOutValid_16 ),
       .io_fabOutValid_15( io_fabOutValid_15 ),
       .io_fabOutValid_14( io_fabOutValid_14 ),
       .io_fabOutValid_13( io_fabOutValid_13 ),
       .io_fabOutValid_12( io_fabOutValid_12 ),
       .io_fabOutValid_11( io_fabOutValid_11 ),
       .io_fabOutValid_10( io_fabOutValid_10 ),
       .io_fabOutValid_9( io_fabOutValid_9 ),
       .io_fabOutValid_8( io_fabOutValid_8 ),
       .io_fabOutValid_7( io_fabOutValid_7 ),
       .io_fabOutValid_6( io_fabOutValid_6 ),
       .io_fabOutValid_5( io_fabOutValid_5 ),
       .io_fabOutValid_4( io_fabOutValid_4 ),
       .io_fabOutValid_3( io_fabOutValid_3 ),
       .io_fabOutValid_2( io_fabOutValid_2 ),
       .io_fabOutValid_1( io_fabOutValid_1 ),
       .io_fabOutValid_0( io_fabOutValid_0 ),
       .io_fabOutRdy_19( fabOutSeqIntClass_io_fabOutRdy_19 ),
       .io_fabOutRdy_18( fabOutSeqIntClass_io_fabOutRdy_18 ),
       .io_fabOutRdy_17( fabOutSeqIntClass_io_fabOutRdy_17 ),
       .io_fabOutRdy_16( fabOutSeqIntClass_io_fabOutRdy_16 ),
       .io_fabOutRdy_15( fabOutSeqIntClass_io_fabOutRdy_15 ),
       .io_fabOutRdy_14( fabOutSeqIntClass_io_fabOutRdy_14 ),
       .io_fabOutRdy_13( fabOutSeqIntClass_io_fabOutRdy_13 ),
       .io_fabOutRdy_12( fabOutSeqIntClass_io_fabOutRdy_12 ),
       .io_fabOutRdy_11( fabOutSeqIntClass_io_fabOutRdy_11 ),
       .io_fabOutRdy_10( fabOutSeqIntClass_io_fabOutRdy_10 ),
       .io_fabOutRdy_9( fabOutSeqIntClass_io_fabOutRdy_9 ),
       .io_fabOutRdy_8( fabOutSeqIntClass_io_fabOutRdy_8 ),
       .io_fabOutRdy_7( fabOutSeqIntClass_io_fabOutRdy_7 ),
       .io_fabOutRdy_6( fabOutSeqIntClass_io_fabOutRdy_6 ),
       .io_fabOutRdy_5( fabOutSeqIntClass_io_fabOutRdy_5 ),
       .io_fabOutRdy_4( fabOutSeqIntClass_io_fabOutRdy_4 ),
       .io_fabOutRdy_3( fabOutSeqIntClass_io_fabOutRdy_3 ),
       .io_fabOutRdy_2( fabOutSeqIntClass_io_fabOutRdy_2 ),
       .io_fabOutRdy_1( fabOutSeqIntClass_io_fabOutRdy_1 ),
       .io_fabOutRdy_0( fabOutSeqIntClass_io_fabOutRdy_0 ),
       .io_fabOutStore_19( fabOutSeqIntClass_io_fabOutStore_19 ),
       .io_fabOutStore_18( fabOutSeqIntClass_io_fabOutStore_18 ),
       .io_fabOutStore_17( fabOutSeqIntClass_io_fabOutStore_17 ),
       .io_fabOutStore_16( fabOutSeqIntClass_io_fabOutStore_16 ),
       .io_fabOutStore_15( fabOutSeqIntClass_io_fabOutStore_15 ),
       .io_fabOutStore_14( fabOutSeqIntClass_io_fabOutStore_14 ),
       .io_fabOutStore_13( fabOutSeqIntClass_io_fabOutStore_13 ),
       .io_fabOutStore_12( fabOutSeqIntClass_io_fabOutStore_12 ),
       .io_fabOutStore_11( fabOutSeqIntClass_io_fabOutStore_11 ),
       .io_fabOutStore_10( fabOutSeqIntClass_io_fabOutStore_10 ),
       .io_fabOutStore_9( fabOutSeqIntClass_io_fabOutStore_9 ),
       .io_fabOutStore_8( fabOutSeqIntClass_io_fabOutStore_8 ),
       .io_fabOutStore_7( fabOutSeqIntClass_io_fabOutStore_7 ),
       .io_fabOutStore_6( fabOutSeqIntClass_io_fabOutStore_6 ),
       .io_fabOutStore_5( fabOutSeqIntClass_io_fabOutStore_5 ),
       .io_fabOutStore_4( fabOutSeqIntClass_io_fabOutStore_4 ),
       .io_fabOutStore_3( fabOutSeqIntClass_io_fabOutStore_3 ),
       .io_fabOutStore_2( fabOutSeqIntClass_io_fabOutStore_2 ),
       .io_fabOutStore_1( fabOutSeqIntClass_io_fabOutStore_1 ),
       .io_fabOutStore_0( fabOutSeqIntClass_io_fabOutStore_0 ),
       .io_fabOutStoreValid_19( fabOutSeqIntClass_io_fabOutStoreValid_19 ),
       .io_fabOutStoreValid_18( fabOutSeqIntClass_io_fabOutStoreValid_18 ),
       .io_fabOutStoreValid_17( fabOutSeqIntClass_io_fabOutStoreValid_17 ),
       .io_fabOutStoreValid_16( fabOutSeqIntClass_io_fabOutStoreValid_16 ),
       .io_fabOutStoreValid_15( fabOutSeqIntClass_io_fabOutStoreValid_15 ),
       .io_fabOutStoreValid_14( fabOutSeqIntClass_io_fabOutStoreValid_14 ),
       .io_fabOutStoreValid_13( fabOutSeqIntClass_io_fabOutStoreValid_13 ),
       .io_fabOutStoreValid_12( fabOutSeqIntClass_io_fabOutStoreValid_12 ),
       .io_fabOutStoreValid_11( fabOutSeqIntClass_io_fabOutStoreValid_11 ),
       .io_fabOutStoreValid_10( fabOutSeqIntClass_io_fabOutStoreValid_10 ),
       .io_fabOutStoreValid_9( fabOutSeqIntClass_io_fabOutStoreValid_9 ),
       .io_fabOutStoreValid_8( fabOutSeqIntClass_io_fabOutStoreValid_8 ),
       .io_fabOutStoreValid_7( fabOutSeqIntClass_io_fabOutStoreValid_7 ),
       .io_fabOutStoreValid_6( fabOutSeqIntClass_io_fabOutStoreValid_6 ),
       .io_fabOutStoreValid_5( fabOutSeqIntClass_io_fabOutStoreValid_5 ),
       .io_fabOutStoreValid_4( fabOutSeqIntClass_io_fabOutStoreValid_4 ),
       .io_fabOutStoreValid_3( fabOutSeqIntClass_io_fabOutStoreValid_3 ),
       .io_fabOutStoreValid_2( fabOutSeqIntClass_io_fabOutStoreValid_2 ),
       .io_fabOutStoreValid_1( fabOutSeqIntClass_io_fabOutStoreValid_1 ),
       .io_fabOutStoreValid_0( fabOutSeqIntClass_io_fabOutStoreValid_0 ),
       .io_fabOutStoreRdy_19( io_fabOutStoreRdy_19 ),
       .io_fabOutStoreRdy_18( io_fabOutStoreRdy_18 ),
       .io_fabOutStoreRdy_17( io_fabOutStoreRdy_17 ),
       .io_fabOutStoreRdy_16( io_fabOutStoreRdy_16 ),
       .io_fabOutStoreRdy_15( io_fabOutStoreRdy_15 ),
       .io_fabOutStoreRdy_14( io_fabOutStoreRdy_14 ),
       .io_fabOutStoreRdy_13( io_fabOutStoreRdy_13 ),
       .io_fabOutStoreRdy_12( io_fabOutStoreRdy_12 ),
       .io_fabOutStoreRdy_11( io_fabOutStoreRdy_11 ),
       .io_fabOutStoreRdy_10( io_fabOutStoreRdy_10 ),
       .io_fabOutStoreRdy_9( io_fabOutStoreRdy_9 ),
       .io_fabOutStoreRdy_8( io_fabOutStoreRdy_8 ),
       .io_fabOutStoreRdy_7( io_fabOutStoreRdy_7 ),
       .io_fabOutStoreRdy_6( io_fabOutStoreRdy_6 ),
       .io_fabOutStoreRdy_5( io_fabOutStoreRdy_5 ),
       .io_fabOutStoreRdy_4( io_fabOutStoreRdy_4 ),
       .io_fabOutStoreRdy_3( io_fabOutStoreRdy_3 ),
       .io_fabOutStoreRdy_2( io_fabOutStoreRdy_2 ),
       .io_fabOutStoreRdy_1( io_fabOutStoreRdy_1 ),
       .io_fabOutStoreRdy_0( io_fabOutStoreRdy_0 ),
       .io_fabOutLoc_19( fabOutSeqIntClass_io_fabOutLoc_19 ),
       .io_fabOutLoc_18( fabOutSeqIntClass_io_fabOutLoc_18 ),
       .io_fabOutLoc_17( fabOutSeqIntClass_io_fabOutLoc_17 ),
       .io_fabOutLoc_16( fabOutSeqIntClass_io_fabOutLoc_16 ),
       .io_fabOutLoc_15( fabOutSeqIntClass_io_fabOutLoc_15 ),
       .io_fabOutLoc_14( fabOutSeqIntClass_io_fabOutLoc_14 ),
       .io_fabOutLoc_13( fabOutSeqIntClass_io_fabOutLoc_13 ),
       .io_fabOutLoc_12( fabOutSeqIntClass_io_fabOutLoc_12 ),
       .io_fabOutLoc_11( fabOutSeqIntClass_io_fabOutLoc_11 ),
       .io_fabOutLoc_10( fabOutSeqIntClass_io_fabOutLoc_10 ),
       .io_fabOutLoc_9( fabOutSeqIntClass_io_fabOutLoc_9 ),
       .io_fabOutLoc_8( fabOutSeqIntClass_io_fabOutLoc_8 ),
       .io_fabOutLoc_7( fabOutSeqIntClass_io_fabOutLoc_7 ),
       .io_fabOutLoc_6( fabOutSeqIntClass_io_fabOutLoc_6 ),
       .io_fabOutLoc_5( fabOutSeqIntClass_io_fabOutLoc_5 ),
       .io_fabOutLoc_4( fabOutSeqIntClass_io_fabOutLoc_4 ),
       .io_fabOutLoc_3( fabOutSeqIntClass_io_fabOutLoc_3 ),
       .io_fabOutLoc_2( fabOutSeqIntClass_io_fabOutLoc_2 ),
       .io_fabOutLoc_1( fabOutSeqIntClass_io_fabOutLoc_1 ),
       .io_fabOutLoc_0( fabOutSeqIntClass_io_fabOutLoc_0 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       .io_fabOutLocRdy_19( fabOutSeqArb_7_io_fabOutLocRdy_19 ),
       .io_fabOutLocRdy_18( fabOutSeqArb_7_io_fabOutLocRdy_18 ),
       .io_fabOutLocRdy_17( fabOutSeqArb_7_io_fabOutLocRdy_17 ),
       .io_fabOutLocRdy_16( fabOutSeqArb_7_io_fabOutLocRdy_16 ),
       .io_fabOutLocRdy_15( fabOutSeqArb_7_io_fabOutLocRdy_15 ),
       .io_fabOutLocRdy_14( fabOutSeqArb_7_io_fabOutLocRdy_14 ),
       .io_fabOutLocRdy_13( fabOutSeqArb_7_io_fabOutLocRdy_13 ),
       .io_fabOutLocRdy_12( fabOutSeqArb_7_io_fabOutLocRdy_12 ),
       .io_fabOutLocRdy_11( fabOutSeqArb_7_io_fabOutLocRdy_11 ),
       .io_fabOutLocRdy_10( fabOutSeqArb_7_io_fabOutLocRdy_10 ),
       .io_fabOutLocRdy_9( fabOutSeqArb_7_io_fabOutLocRdy_9 ),
       .io_fabOutLocRdy_8( fabOutSeqArb_7_io_fabOutLocRdy_8 ),
       .io_fabOutLocRdy_7( fabOutSeqArb_7_io_fabOutLocRdy_7 ),
       .io_fabOutLocRdy_6( fabOutSeqArb_7_io_fabOutLocRdy_6 ),
       .io_fabOutLocRdy_5( fabOutSeqArb_7_io_fabOutLocRdy_5 ),
       .io_fabOutLocRdy_4( fabOutSeqArb_7_io_fabOutLocRdy_4 ),
       .io_fabOutLocRdy_3( fabOutSeqArb_7_io_fabOutLocRdy_3 ),
       .io_fabOutLocRdy_2( fabOutSeqArb_7_io_fabOutLocRdy_2 ),
       .io_fabOutLocRdy_1( fabOutSeqArb_7_io_fabOutLocRdy_1 ),
       .io_fabOutLocRdy_0( fabOutSeqArb_7_io_fabOutLocRdy_0 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T159 ),
       .io_fabOutLoc_18( T158 ),
       .io_fabOutLoc_17( T157 ),
       .io_fabOutLoc_16( T156 ),
       .io_fabOutLoc_15( T155 ),
       .io_fabOutLoc_14( T154 ),
       .io_fabOutLoc_13( T153 ),
       .io_fabOutLoc_12( T152 ),
       .io_fabOutLoc_11( T151 ),
       .io_fabOutLoc_10( T150 ),
       .io_fabOutLoc_9( T149 ),
       .io_fabOutLoc_8( T148 ),
       .io_fabOutLoc_7( T147 ),
       .io_fabOutLoc_6( T146 ),
       .io_fabOutLoc_5( T145 ),
       .io_fabOutLoc_4( T144 ),
       .io_fabOutLoc_3( T143 ),
       .io_fabOutLoc_2( T142 ),
       .io_fabOutLoc_1( T141 ),
       .io_fabOutLoc_0( T140 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_0 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_1(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T139 ),
       .io_fabOutLoc_18( T138 ),
       .io_fabOutLoc_17( T137 ),
       .io_fabOutLoc_16( T136 ),
       .io_fabOutLoc_15( T135 ),
       .io_fabOutLoc_14( T134 ),
       .io_fabOutLoc_13( T133 ),
       .io_fabOutLoc_12( T132 ),
       .io_fabOutLoc_11( T131 ),
       .io_fabOutLoc_10( T130 ),
       .io_fabOutLoc_9( T129 ),
       .io_fabOutLoc_8( T128 ),
       .io_fabOutLoc_7( T127 ),
       .io_fabOutLoc_6( T126 ),
       .io_fabOutLoc_5( T125 ),
       .io_fabOutLoc_4( T124 ),
       .io_fabOutLoc_3( T123 ),
       .io_fabOutLoc_2( T122 ),
       .io_fabOutLoc_1( T121 ),
       .io_fabOutLoc_0( T120 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_1_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_1_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_1 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_2(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T119 ),
       .io_fabOutLoc_18( T118 ),
       .io_fabOutLoc_17( T117 ),
       .io_fabOutLoc_16( T116 ),
       .io_fabOutLoc_15( T115 ),
       .io_fabOutLoc_14( T114 ),
       .io_fabOutLoc_13( T113 ),
       .io_fabOutLoc_12( T112 ),
       .io_fabOutLoc_11( T111 ),
       .io_fabOutLoc_10( T110 ),
       .io_fabOutLoc_9( T109 ),
       .io_fabOutLoc_8( T108 ),
       .io_fabOutLoc_7( T107 ),
       .io_fabOutLoc_6( T106 ),
       .io_fabOutLoc_5( T105 ),
       .io_fabOutLoc_4( T104 ),
       .io_fabOutLoc_3( T103 ),
       .io_fabOutLoc_2( T102 ),
       .io_fabOutLoc_1( T101 ),
       .io_fabOutLoc_0( T100 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_2_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_2_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_2 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_3(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T99 ),
       .io_fabOutLoc_18( T98 ),
       .io_fabOutLoc_17( T97 ),
       .io_fabOutLoc_16( T96 ),
       .io_fabOutLoc_15( T95 ),
       .io_fabOutLoc_14( T94 ),
       .io_fabOutLoc_13( T93 ),
       .io_fabOutLoc_12( T92 ),
       .io_fabOutLoc_11( T91 ),
       .io_fabOutLoc_10( T90 ),
       .io_fabOutLoc_9( T89 ),
       .io_fabOutLoc_8( T88 ),
       .io_fabOutLoc_7( T87 ),
       .io_fabOutLoc_6( T86 ),
       .io_fabOutLoc_5( T85 ),
       .io_fabOutLoc_4( T84 ),
       .io_fabOutLoc_3( T83 ),
       .io_fabOutLoc_2( T82 ),
       .io_fabOutLoc_1( T81 ),
       .io_fabOutLoc_0( T80 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_3_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_3_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_3 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_4(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T79 ),
       .io_fabOutLoc_18( T78 ),
       .io_fabOutLoc_17( T77 ),
       .io_fabOutLoc_16( T76 ),
       .io_fabOutLoc_15( T75 ),
       .io_fabOutLoc_14( T74 ),
       .io_fabOutLoc_13( T73 ),
       .io_fabOutLoc_12( T72 ),
       .io_fabOutLoc_11( T71 ),
       .io_fabOutLoc_10( T70 ),
       .io_fabOutLoc_9( T69 ),
       .io_fabOutLoc_8( T68 ),
       .io_fabOutLoc_7( T67 ),
       .io_fabOutLoc_6( T66 ),
       .io_fabOutLoc_5( T65 ),
       .io_fabOutLoc_4( T64 ),
       .io_fabOutLoc_3( T63 ),
       .io_fabOutLoc_2( T62 ),
       .io_fabOutLoc_1( T61 ),
       .io_fabOutLoc_0( T60 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_4_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_4_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_4 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_5(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T59 ),
       .io_fabOutLoc_18( T58 ),
       .io_fabOutLoc_17( T57 ),
       .io_fabOutLoc_16( T56 ),
       .io_fabOutLoc_15( T55 ),
       .io_fabOutLoc_14( T54 ),
       .io_fabOutLoc_13( T53 ),
       .io_fabOutLoc_12( T52 ),
       .io_fabOutLoc_11( T51 ),
       .io_fabOutLoc_10( T50 ),
       .io_fabOutLoc_9( T49 ),
       .io_fabOutLoc_8( T48 ),
       .io_fabOutLoc_7( T47 ),
       .io_fabOutLoc_6( T46 ),
       .io_fabOutLoc_5( T45 ),
       .io_fabOutLoc_4( T44 ),
       .io_fabOutLoc_3( T43 ),
       .io_fabOutLoc_2( T42 ),
       .io_fabOutLoc_1( T41 ),
       .io_fabOutLoc_0( T40 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_5_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_5_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_5 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_6(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T39 ),
       .io_fabOutLoc_18( T38 ),
       .io_fabOutLoc_17( T37 ),
       .io_fabOutLoc_16( T36 ),
       .io_fabOutLoc_15( T35 ),
       .io_fabOutLoc_14( T34 ),
       .io_fabOutLoc_13( T33 ),
       .io_fabOutLoc_12( T32 ),
       .io_fabOutLoc_11( T31 ),
       .io_fabOutLoc_10( T30 ),
       .io_fabOutLoc_9( T29 ),
       .io_fabOutLoc_8( T28 ),
       .io_fabOutLoc_7( T27 ),
       .io_fabOutLoc_6( T26 ),
       .io_fabOutLoc_5( T25 ),
       .io_fabOutLoc_4( T24 ),
       .io_fabOutLoc_3( T23 ),
       .io_fabOutLoc_2( T22 ),
       .io_fabOutLoc_1( T21 ),
       .io_fabOutLoc_0( T20 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       //.io_fabOutLocRdy_19(  )
       //.io_fabOutLocRdy_18(  )
       //.io_fabOutLocRdy_17(  )
       //.io_fabOutLocRdy_16(  )
       //.io_fabOutLocRdy_15(  )
       //.io_fabOutLocRdy_14(  )
       //.io_fabOutLocRdy_13(  )
       //.io_fabOutLocRdy_12(  )
       //.io_fabOutLocRdy_11(  )
       //.io_fabOutLocRdy_10(  )
       //.io_fabOutLocRdy_9(  )
       //.io_fabOutLocRdy_8(  )
       //.io_fabOutLocRdy_7(  )
       //.io_fabOutLocRdy_6(  )
       //.io_fabOutLocRdy_5(  )
       //.io_fabOutLocRdy_4(  )
       //.io_fabOutLocRdy_3(  )
       //.io_fabOutLocRdy_2(  )
       //.io_fabOutLocRdy_1(  )
       //.io_fabOutLocRdy_0(  )
       .io_locStoreData( fabOutSeqArb_6_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_6_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_6 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
  fabOutSeqArb fabOutSeqArb_7(.clk(clk), .reset(reset),
       .io_fabOutLoc_19( T19 ),
       .io_fabOutLoc_18( T18 ),
       .io_fabOutLoc_17( T17 ),
       .io_fabOutLoc_16( T16 ),
       .io_fabOutLoc_15( T15 ),
       .io_fabOutLoc_14( T14 ),
       .io_fabOutLoc_13( T13 ),
       .io_fabOutLoc_12( T12 ),
       .io_fabOutLoc_11( T11 ),
       .io_fabOutLoc_10( T10 ),
       .io_fabOutLoc_9( T9 ),
       .io_fabOutLoc_8( T8 ),
       .io_fabOutLoc_7( T7 ),
       .io_fabOutLoc_6( T6 ),
       .io_fabOutLoc_5( T5 ),
       .io_fabOutLoc_4( T4 ),
       .io_fabOutLoc_3( T3 ),
       .io_fabOutLoc_2( T2 ),
       .io_fabOutLoc_1( T1 ),
       .io_fabOutLoc_0( T0 ),
       .io_fabOutLocValid_19( fabOutSeqIntClass_io_fabOutLocValid_19 ),
       .io_fabOutLocValid_18( fabOutSeqIntClass_io_fabOutLocValid_18 ),
       .io_fabOutLocValid_17( fabOutSeqIntClass_io_fabOutLocValid_17 ),
       .io_fabOutLocValid_16( fabOutSeqIntClass_io_fabOutLocValid_16 ),
       .io_fabOutLocValid_15( fabOutSeqIntClass_io_fabOutLocValid_15 ),
       .io_fabOutLocValid_14( fabOutSeqIntClass_io_fabOutLocValid_14 ),
       .io_fabOutLocValid_13( fabOutSeqIntClass_io_fabOutLocValid_13 ),
       .io_fabOutLocValid_12( fabOutSeqIntClass_io_fabOutLocValid_12 ),
       .io_fabOutLocValid_11( fabOutSeqIntClass_io_fabOutLocValid_11 ),
       .io_fabOutLocValid_10( fabOutSeqIntClass_io_fabOutLocValid_10 ),
       .io_fabOutLocValid_9( fabOutSeqIntClass_io_fabOutLocValid_9 ),
       .io_fabOutLocValid_8( fabOutSeqIntClass_io_fabOutLocValid_8 ),
       .io_fabOutLocValid_7( fabOutSeqIntClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqIntClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqIntClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqIntClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqIntClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqIntClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqIntClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqIntClass_io_fabOutLocValid_0 ),
       .io_fabOutLocRdy_19( fabOutSeqArb_7_io_fabOutLocRdy_19 ),
       .io_fabOutLocRdy_18( fabOutSeqArb_7_io_fabOutLocRdy_18 ),
       .io_fabOutLocRdy_17( fabOutSeqArb_7_io_fabOutLocRdy_17 ),
       .io_fabOutLocRdy_16( fabOutSeqArb_7_io_fabOutLocRdy_16 ),
       .io_fabOutLocRdy_15( fabOutSeqArb_7_io_fabOutLocRdy_15 ),
       .io_fabOutLocRdy_14( fabOutSeqArb_7_io_fabOutLocRdy_14 ),
       .io_fabOutLocRdy_13( fabOutSeqArb_7_io_fabOutLocRdy_13 ),
       .io_fabOutLocRdy_12( fabOutSeqArb_7_io_fabOutLocRdy_12 ),
       .io_fabOutLocRdy_11( fabOutSeqArb_7_io_fabOutLocRdy_11 ),
       .io_fabOutLocRdy_10( fabOutSeqArb_7_io_fabOutLocRdy_10 ),
       .io_fabOutLocRdy_9( fabOutSeqArb_7_io_fabOutLocRdy_9 ),
       .io_fabOutLocRdy_8( fabOutSeqArb_7_io_fabOutLocRdy_8 ),
       .io_fabOutLocRdy_7( fabOutSeqArb_7_io_fabOutLocRdy_7 ),
       .io_fabOutLocRdy_6( fabOutSeqArb_7_io_fabOutLocRdy_6 ),
       .io_fabOutLocRdy_5( fabOutSeqArb_7_io_fabOutLocRdy_5 ),
       .io_fabOutLocRdy_4( fabOutSeqArb_7_io_fabOutLocRdy_4 ),
       .io_fabOutLocRdy_3( fabOutSeqArb_7_io_fabOutLocRdy_3 ),
       .io_fabOutLocRdy_2( fabOutSeqArb_7_io_fabOutLocRdy_2 ),
       .io_fabOutLocRdy_1( fabOutSeqArb_7_io_fabOutLocRdy_1 ),
       .io_fabOutLocRdy_0( fabOutSeqArb_7_io_fabOutLocRdy_0 ),
       .io_locStoreData( fabOutSeqArb_7_io_locStoreData ),
       .io_locStoreValid( fabOutSeqArb_7_io_locStoreValid ),
       .io_locStoreRdy( io_fabOutLocRdy_7 ),
       .io_rst( fabOutSeqIntClass_io_rst )
  );
endmodule

module controllerConfigure_1(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_outConfig,
    output io_outValid,
    output io_computeCtrl,
    output io_computeCtrlValid
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  reg [31:0] inDataReg;
  wire[31:0] T30;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inDataReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_computeCtrlValid = T0;
  assign T0 = T21 ? 1'h0 : T1;
  assign T1 = T18 ? 1'h1 : T2;
  assign T2 = T13 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : 1'h0;
  assign T4 = T11 & T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 2'h0;
  assign T7 = inDataReg[5'h1f:5'h1e];
  assign T30 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inDataReg;
  assign T9 = T10 == 1'h1;
  assign T10 = inDataReg[1'h0:1'h0];
  assign T11 = T12 == 1'h0;
  assign T12 = inDataReg[5'h1f:5'h1f];
  assign T13 = T11 & T14;
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inDataReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T11 & T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T5 | T15;
  assign T21 = T11 ^ 1'h1;
  assign io_computeCtrl = T22;
  assign T22 = T21 ? 1'h0 : T23;
  assign T23 = T18 ? 1'h0 : T24;
  assign T24 = T13 ? 1'h0 : T25;
  assign T25 = T4 ? 1'h1 : 1'h0;
  assign io_outValid = T26;
  assign T26 = T21 ? 1'h0 : T27;
  assign T27 = T18 ? 1'h0 : T28;
  assign T28 = T13 ? 1'h1 : T29;
  assign T29 = T4 ? 1'h0 : 1'h0;
  assign io_outConfig = inDataReg;

  always @(posedge clk) begin
    if(reset) begin
      inDataReg <= 32'h0;
    end else if(io_inValid) begin
      inDataReg <= io_inConfig;
    end
  end
endmodule

module loadSeqCtrl(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output io_spillEnd,
    output io_nextIterStart,
    output[8:0] io_seqMemAddr,
    output io_seqMemAddrValid,
    output io_computeEnable,
    input  io_seqProceed
);

  reg  computeEnable;
  wire T124;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[514:0] lastAddr;
  wire[514:0] T125;
  wire[513:0] T6;
  wire[513:0] T126;
  reg [8:0] epilogueDepth;
  wire[8:0] T127;
  wire[8:0] T7;
  wire[8:0] T128;
  wire[6:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[9:0] T21;
  wire[513:0] ssEnd;
  wire[513:0] T129;
  wire[8:0] T22;
  reg [8:0] steadyStateDepth;
  wire[8:0] T130;
  wire[9:0] T131;
  wire[9:0] T23;
  wire[9:0] T132;
  wire[9:0] T24;
  wire T25;
  reg [8:0] prologueDepth;
  wire[8:0] T133;
  wire[8:0] T26;
  wire[8:0] T134;
  wire[6:0] T27;
  wire startComputeValid;
  wire T28;
  wire T29;
  wire computeCtrl;
  wire computeCtrlValid;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire computeDone;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[514:0] T39;
  wire[514:0] T135;
  reg [511:0] seqMemAddr;
  wire[511:0] T136;
  wire[513:0] T137;
  wire[513:0] T40;
  wire[513:0] T41;
  wire[513:0] T138;
  wire[511:0] T42;
  wire[511:0] T43;
  wire[511:0] T44;
  wire T45;
  wire T46;
  wire nextRequest;
  wire[511:0] T139;
  wire T47;
  wire T48;
  wire T49;
  reg [8:0] epilogueSpill;
  wire[8:0] T140;
  wire[9:0] T141;
  wire[9:0] T50;
  wire[9:0] T142;
  wire[9:0] T51;
  wire T52;
  wire[31:0] T53;
  reg [31:0] iterCount;
  wire[31:0] T143;
  wire[31:0] T54;
  wire[31:0] T144;
  wire[18:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[2:0] T59;
  wire T60;
  reg [31:0] currentIter;
  wire[31:0] T145;
  wire[31:0] T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire T64;
  wire T65;
  wire[513:0] T66;
  wire[513:0] T146;
  wire T67;
  wire T68;
  wire[511:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[511:0] T147;
  wire T76;
  reg  spillEnd;
  wire T148;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[513:0] T149;
  wire[511:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire[514:0] T96;
  wire[514:0] T150;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[513:0] T104;
  wire[513:0] spillEndAddr;
  wire[513:0] T151;
  wire[8:0] T105;
  wire[513:0] T152;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire resetComputeValid;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[8:0] T153;
  reg  nextIterStart;
  wire T154;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire loadCtrlConfigure_io_computeCtrl;
  wire loadCtrlConfigure_io_computeCtrlValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    computeEnable = {1{$random}};
    epilogueDepth = {1{$random}};
    steadyStateDepth = {1{$random}};
    prologueDepth = {1{$random}};
    seqMemAddr = {16{$random}};
    epilogueSpill = {1{$random}};
    iterCount = {1{$random}};
    currentIter = {1{$random}};
    spillEnd = {1{$random}};
    nextIterStart = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign io_seqMemAddrValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_computeEnable = computeEnable;
  assign T124 = reset ? 1'h0 : T0;
  assign T0 = T116 ? 1'h0 : T1;
  assign T1 = T113 ? 1'h0 : T2;
  assign T2 = T3 ? 1'h1 : computeEnable;
  assign T3 = T34 & T4;
  assign T4 = startComputeValid & T5;
  assign T5 = lastAddr != 515'h0;
  assign lastAddr = T125;
  assign T125 = {1'h0, T6};
  assign T6 = ssEnd + T126;
  assign T126 = {505'h0, epilogueDepth};
  assign T127 = reset ? 9'h0 : T7;
  assign T7 = T9 ? T128 : epilogueDepth;
  assign T128 = {2'h0, T8};
  assign T8 = io_inConfig[3'h6:1'h0];
  assign T9 = T16 & T10;
  assign T10 = T13 & T11;
  assign T11 = T12 == 1'h1;
  assign T12 = io_inConfig[5'h11:5'h11];
  assign T13 = T14 ^ 1'h1;
  assign T14 = T15 == 1'h0;
  assign T15 = io_inConfig[5'h11:5'h11];
  assign T16 = T19 & T17;
  assign T17 = T18 == 3'h0;
  assign T18 = io_inConfig[5'h15:5'h13];
  assign T19 = io_inValid & T20;
  assign T20 = T21 == 10'h100;
  assign T21 = io_inConfig[5'h1f:5'h16];
  assign ssEnd = T129;
  assign T129 = {505'h0, T22};
  assign T22 = prologueDepth + steadyStateDepth;
  assign T130 = T131[4'h8:1'h0];
  assign T131 = reset ? 10'h0 : T23;
  assign T23 = T25 ? T24 : T132;
  assign T132 = {1'h0, steadyStateDepth};
  assign T24 = io_inConfig[5'h10:3'h7];
  assign T25 = T16 & T14;
  assign T133 = reset ? 9'h0 : T26;
  assign T26 = T25 ? T134 : prologueDepth;
  assign T134 = {2'h0, T27};
  assign T27 = io_inConfig[3'h6:1'h0];
  assign startComputeValid = T28;
  assign T28 = T30 ? 1'h0 : T29;
  assign T29 = computeCtrlValid & computeCtrl;
  assign computeCtrl = loadCtrlConfigure_io_computeCtrl;
  assign computeCtrlValid = loadCtrlConfigure_io_computeCtrlValid;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T29 | T32;
  assign T32 = computeCtrlValid & T33;
  assign T33 = computeCtrl ^ 1'h1;
  assign T34 = T109 | computeDone;
  assign computeDone = T35;
  assign T35 = T106 ? T101 : T36;
  assign T36 = T97 ? T92 : T37;
  assign T37 = T87 ? T38 : 1'h0;
  assign T38 = T135 == T39;
  assign T39 = lastAddr - 515'h1;
  assign T135 = {3'h0, seqMemAddr};
  assign T136 = T137[9'h1ff:1'h0];
  assign T137 = reset ? 514'h0 : T40;
  assign T40 = T84 ? T149 : T41;
  assign T41 = T72 ? ssEnd : T138;
  assign T138 = {2'h0, T42};
  assign T42 = T70 ? T69 : T43;
  assign T43 = T47 ? T139 : T44;
  assign T44 = T45 ? 512'h0 : seqMemAddr;
  assign T45 = T46 & startComputeValid;
  assign T46 = startComputeValid | nextRequest;
  assign nextRequest = io_seqProceed;
  assign T139 = {503'h0, prologueDepth};
  assign T47 = T64 & T48;
  assign T48 = T52 | T49;
  assign T49 = epilogueSpill != 9'h0;
  assign T140 = T141[4'h8:1'h0];
  assign T141 = reset ? 10'h0 : T50;
  assign T50 = T9 ? T51 : T142;
  assign T142 = {1'h0, epilogueSpill};
  assign T51 = io_inConfig[5'h10:3'h7];
  assign T52 = currentIter < T53;
  assign T53 = iterCount - 32'h1;
  assign T143 = reset ? 32'h0 : T54;
  assign T54 = T56 ? T144 : iterCount;
  assign T144 = {13'h0, T55};
  assign T55 = io_inConfig[5'h12:1'h0];
  assign T56 = T19 & T57;
  assign T57 = T60 & T58;
  assign T58 = T59 == 3'h0;
  assign T59 = io_inConfig[5'h15:5'h13];
  assign T60 = T17 ^ 1'h1;
  assign T145 = reset ? 32'h0 : T61;
  assign T61 = T47 ? T63 : T62;
  assign T62 = T45 ? 32'h0 : currentIter;
  assign T63 = currentIter + 32'h1;
  assign T64 = T67 & T65;
  assign T65 = T146 == T66;
  assign T66 = ssEnd - 514'h1;
  assign T146 = {2'h0, seqMemAddr};
  assign T67 = T46 & T68;
  assign T68 = startComputeValid ^ 1'h1;
  assign T69 = seqMemAddr + 512'h1;
  assign T70 = T64 & T71;
  assign T71 = T48 ^ 1'h1;
  assign T72 = T67 & T73;
  assign T73 = T82 & T74;
  assign T74 = T81 & T75;
  assign T75 = seqMemAddr == T147;
  assign T147 = {511'h0, T76};
  assign T76 = spillEnd - 1'h1;
  assign T148 = reset ? 1'h0 : T77;
  assign T77 = T84 ? 1'h0 : T78;
  assign T78 = T72 ? 1'h1 : T79;
  assign T79 = T64 ? 1'h0 : T80;
  assign T80 = T45 ? 1'h0 : spillEnd;
  assign T81 = currentIter == iterCount;
  assign T82 = T65 ^ 1'h1;
  assign T149 = {2'h0, T83};
  assign T83 = seqMemAddr + 512'h1;
  assign T84 = T67 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T65 | T74;
  assign T87 = T91 & T88;
  assign T88 = T90 & T89;
  assign T89 = steadyStateDepth == 9'h0;
  assign T90 = epilogueDepth != 9'h0;
  assign T91 = computeEnable & nextRequest;
  assign T92 = T95 & T93;
  assign T93 = T94 == iterCount;
  assign T94 = currentIter + 32'h1;
  assign T95 = T150 == T96;
  assign T96 = lastAddr - 515'h1;
  assign T150 = {3'h0, seqMemAddr};
  assign T97 = T91 & T98;
  assign T98 = T100 & T99;
  assign T99 = epilogueSpill == 9'h0;
  assign T100 = T88 ^ 1'h1;
  assign T101 = T103 & T102;
  assign T102 = currentIter == iterCount;
  assign T103 = T152 == T104;
  assign T104 = spillEndAddr - 514'h1;
  assign spillEndAddr = T151;
  assign T151 = {505'h0, T105};
  assign T105 = prologueDepth + epilogueSpill;
  assign T152 = {2'h0, seqMemAddr};
  assign T106 = T91 & T107;
  assign T107 = T108 ^ 1'h1;
  assign T108 = T88 | T99;
  assign T109 = startComputeValid | resetComputeValid;
  assign resetComputeValid = T110;
  assign T110 = T30 ? 1'h0 : T111;
  assign T111 = T112 & T32;
  assign T112 = T29 ^ 1'h1;
  assign T113 = T34 & T114;
  assign T114 = T115 & resetComputeValid;
  assign T115 = T4 ^ 1'h1;
  assign T116 = T34 & T117;
  assign T117 = T118 ^ 1'h1;
  assign T118 = T4 | resetComputeValid;
  assign io_seqMemAddr = T153;
  assign T153 = seqMemAddr[4'h8:1'h0];
  assign io_nextIterStart = nextIterStart;
  assign T154 = reset ? 1'h0 : T119;
  assign T119 = T84 ? 1'h0 : T120;
  assign T120 = T72 ? 1'h0 : T121;
  assign T121 = T70 ? 1'h0 : T122;
  assign T122 = T47 ? 1'h1 : T123;
  assign T123 = T45 ? 1'h0 : nextIterStart;
  assign io_spillEnd = spillEnd;
  controllerConfigure_1 loadCtrlConfigure(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       //.io_outConfig(  )
       //.io_outValid(  )
       .io_computeCtrl( loadCtrlConfigure_io_computeCtrl ),
       .io_computeCtrlValid( loadCtrlConfigure_io_computeCtrlValid )
  );

  always @(posedge clk) begin
    if(reset) begin
      computeEnable <= 1'h0;
    end else if(T116) begin
      computeEnable <= 1'h0;
    end else if(T113) begin
      computeEnable <= 1'h0;
    end else if(T3) begin
      computeEnable <= 1'h1;
    end
    if(reset) begin
      epilogueDepth <= 9'h0;
    end else if(T9) begin
      epilogueDepth <= T128;
    end
    steadyStateDepth <= T130;
    if(reset) begin
      prologueDepth <= 9'h0;
    end else if(T25) begin
      prologueDepth <= T134;
    end
    seqMemAddr <= T136;
    epilogueSpill <= T140;
    if(reset) begin
      iterCount <= 32'h0;
    end else if(T56) begin
      iterCount <= T144;
    end
    if(reset) begin
      currentIter <= 32'h0;
    end else if(T47) begin
      currentIter <= T63;
    end else if(T45) begin
      currentIter <= 32'h0;
    end
    if(reset) begin
      spillEnd <= 1'h0;
    end else if(T84) begin
      spillEnd <= 1'h0;
    end else if(T72) begin
      spillEnd <= 1'h1;
    end else if(T64) begin
      spillEnd <= 1'h0;
    end else if(T45) begin
      spillEnd <= 1'h0;
    end
    if(reset) begin
      nextIterStart <= 1'h0;
    end else if(T84) begin
      nextIterStart <= 1'h0;
    end else if(T72) begin
      nextIterStart <= 1'h0;
    end else if(T70) begin
      nextIterStart <= 1'h0;
    end else if(T47) begin
      nextIterStart <= 1'h1;
    end else if(T45) begin
      nextIterStart <= 1'h0;
    end
  end
endmodule

module customReg_1(input clk,
    input [31:0] io_inData,
    output[31:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [4:0] io_readAddr,
    input [4:0] io_writeAddr
);

  wire[31:0] T0;
  reg [31:0] ram [19:0];
  wire[31:0] T1;
  wire T2;
  wire T3;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 20; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];
  assign T2 = io_writeEn & T3;
  assign T3 = io_writeAddr < 5'h14;

  always @(posedge clk) begin
    if (T2)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module customReg_2(input clk,
    input [56:0] io_inData,
    output[56:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [5:0] io_readAddr,
    input [5:0] io_writeAddr
);

  wire[56:0] T0;
  reg [56:0] ram [59:0];
  wire[56:0] T1;
  wire T2;
  wire T3;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 60; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];
  assign T2 = io_writeEn & T3;
  assign T3 = io_writeAddr < 6'h3c;

  always @(posedge clk) begin
    if (T2)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module customReg_3(input clk,
    input [42:0] io_inData,
    output[42:0] io_outData,
    input  io_readEn,
    input  io_writeEn,
    input [8:0] io_readAddr,
    input [8:0] io_writeAddr
);

  wire[42:0] T0;
  reg [42:0] ram [511:0];
  wire[42:0] T1;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 512; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_outData = T0;
  assign T0 = ram[io_readAddr];

  always @(posedge clk) begin
    if (io_writeEn)
      ram[io_writeAddr] <= io_inData;
  end
endmodule

module memConfig_1(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[8:0] io_memAddr,
    output[42:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[42:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[8:0] T87;
  reg [8:0] memAddr;
  wire[8:0] T97;
  wire[8:0] T88;
  wire[8:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h2;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h2;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h2;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h2;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[6'h2a:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 9'h0;
  assign T97 = reset ? 9'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 9'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 9'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_2(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[5:0] io_memAddr,
    output[56:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[56:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[5:0] T87;
  reg [5:0] memAddr;
  wire[5:0] T97;
  wire[5:0] T88;
  wire[5:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h3;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h3;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h3;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h3;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[6'h38:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 6'h0;
  assign T97 = reset ? 6'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 6'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 6'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_3(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T97;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h4;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h4;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h4;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h4;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T97 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_4(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T97;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h5;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h5;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h5;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h5;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T97 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_5(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T94;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T95;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T96;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T97;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T58 == 5'h6;
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T63 == 5'h6;
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T68 == 5'h6;
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T73 == 5'h6;
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T94;
  assign T94 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T95 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T96 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T97 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module fifo_2(input clk, input reset,
    input [37:0] io_enqData,
    output[37:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg [2:0] deqPtr;
  wire[2:0] T21;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] deqPtrInc;
  wire[2:0] T4;
  wire doDeq;
  wire T5;
  reg [2:0] enqPtr;
  wire[2:0] T22;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] enqPtrInc;
  wire[2:0] T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[37:0] T19;
  reg [37:0] fifoMem [7:0];
  wire[37:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 3'h0 : T2;
  assign T2 = io_rst ? 3'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 4'h8;
  assign T4 = deqPtr + 3'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 3'h0 : T6;
  assign T6 = io_rst ? 3'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 4'h8;
  assign T8 = enqPtr + 3'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 3'h0;
    end else if(io_rst) begin
      deqPtr <= 3'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 3'h0;
    end else if(io_rst) begin
      enqPtr <= 3'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fifo_3(input clk, input reset,
    input [31:0] io_enqData,
    output[31:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg [2:0] deqPtr;
  wire[2:0] T21;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] deqPtrInc;
  wire[2:0] T4;
  wire doDeq;
  wire T5;
  reg [2:0] enqPtr;
  wire[2:0] T22;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] enqPtrInc;
  wire[2:0] T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[31:0] T19;
  reg [31:0] fifoMem [7:0];
  wire[31:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      fifoMem[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 3'h0 : T2;
  assign T2 = io_rst ? 3'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 4'h8;
  assign T4 = deqPtr + 3'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 3'h0 : T6;
  assign T6 = io_rst ? 3'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 4'h8;
  assign T8 = enqPtr + 3'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 3'h0;
    end else if(io_rst) begin
      deqPtr <= 3'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 3'h0;
    end else if(io_rst) begin
      enqPtr <= 3'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module fifo_4(input clk, input reset,
    input [37:0] io_enqData,
    output[37:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg  deqPtr;
  wire T21;
  wire T2;
  wire T3;
  wire deqPtrInc;
  wire T4;
  wire doDeq;
  wire T5;
  reg  enqPtr;
  wire T22;
  wire T6;
  wire T7;
  wire enqPtrInc;
  wire T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[37:0] T19;
  reg [37:0] fifoMem [1:0];
  wire[37:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = io_rst ? 1'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 2'h2;
  assign T4 = deqPtr + 1'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 1'h0 : T6;
  assign T6 = io_rst ? 1'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 2'h2;
  assign T8 = enqPtr + 1'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 1'h0;
    end else if(io_rst) begin
      deqPtr <= 1'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 1'h0;
    end else if(io_rst) begin
      enqPtr <= 1'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module loadSeqDP(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input  io_spillEnd,
    input  io_nextIterStart,
    input [8:0] io_seqMemAddr,
    input  io_seqMemAddrValid,
    output[37:0] io_memBankEnq_7,
    output[37:0] io_memBankEnq_6,
    output[37:0] io_memBankEnq_5,
    output[37:0] io_memBankEnq_4,
    output[37:0] io_memBankEnq_3,
    output[37:0] io_memBankEnq_2,
    output[37:0] io_memBankEnq_1,
    output[37:0] io_memBankEnq_0,
    output io_memBankValid_7,
    output io_memBankValid_6,
    output io_memBankValid_5,
    output io_memBankValid_4,
    output io_memBankValid_3,
    output io_memBankValid_2,
    output io_memBankValid_1,
    output io_memBankValid_0,
    input  io_memBankRdy_7,
    input  io_memBankRdy_6,
    input  io_memBankRdy_5,
    input  io_memBankRdy_4,
    input  io_memBankRdy_3,
    input  io_memBankRdy_2,
    input  io_memBankRdy_1,
    input  io_memBankRdy_0,
    output[31:0] io_loadRqst,
    output io_loadRqstValid,
    input  io_loadRqstRdy,
    input [37:0] io_loadResp,
    input  io_loadRespValid,
    output io_loadRespRdy,
    output io_seqProceed
);

  wire T0;
  wire T1;
  wire T2;
  wire enqReqWire_7;
  wire T3;
  wire T4;
  reg [56:0] lRespDest;
  wire[56:0] T746;
  wire[56:0] T5;
  wire[56:0] regLookup;
  wire[56:0] T6;
  wire T7;
  wire enqComplete;
  wire T8;
  wire T9;
  reg [7:0] enqDoneReg;
  wire[7:0] T747;
  wire[7:0] T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire[7:0] T16;
  wire[7:0] T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T748;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[7:0] T26;
  wire[7:0] T27;
  wire[7:0] T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T749;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire enqReqWire_6;
  wire T36;
  wire T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T750;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire enqReqWire_5;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T751;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire enqReqWire_4;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T752;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire enqReqWire_3;
  wire T72;
  wire T73;
  wire[7:0] T74;
  wire[7:0] T75;
  wire[7:0] T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T753;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire enqReqWire_2;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T754;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire enqReqWire_1;
  wire T96;
  wire T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T755;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire enqReqWire_0;
  wire T108;
  wire T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T756;
  wire T116;
  wire T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T757;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire[7:0] T128;
  wire T129;
  wire[7:0] T130;
  wire[7:0] T131;
  wire[7:0] T132;
  wire[7:0] T133;
  wire[7:0] T758;
  wire T134;
  wire T135;
  wire[7:0] T136;
  wire[7:0] T137;
  wire T138;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[7:0] T141;
  wire[7:0] T142;
  wire[7:0] T759;
  wire T143;
  wire T144;
  wire[7:0] T145;
  wire[7:0] T146;
  wire T147;
  wire[7:0] T148;
  wire[7:0] T149;
  wire[7:0] T150;
  wire[7:0] T151;
  wire[7:0] T760;
  wire T152;
  wire T153;
  wire[7:0] T154;
  wire[7:0] T155;
  wire T156;
  wire[7:0] T157;
  wire[7:0] T158;
  wire[7:0] T159;
  wire[7:0] T160;
  wire[7:0] T761;
  wire T161;
  wire T162;
  wire[7:0] T163;
  wire[7:0] T164;
  wire T165;
  wire[7:0] T166;
  wire[7:0] T167;
  wire[7:0] T168;
  wire[7:0] T169;
  wire[7:0] T762;
  wire T170;
  wire T171;
  wire[7:0] T172;
  wire[7:0] T173;
  wire T174;
  wire[7:0] T175;
  wire[7:0] T176;
  wire[7:0] T177;
  wire[7:0] T178;
  wire[7:0] T763;
  wire T179;
  wire T180;
  wire[7:0] T181;
  wire[7:0] T182;
  reg  lRespLkupValid;
  wire T764;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[37:0] T188;
  wire[37:0] T189;
  wire[31:0] T190;
  reg [31:0] lRespData;
  wire[31:0] T765;
  wire[31:0] T191;
  wire[31:0] regLookupData;
  wire[31:0] T192;
  wire[31:0] T193;
  wire[5:0] T194;
  wire T195;
  wire T196;
  wire[37:0] T197;
  wire[37:0] T198;
  wire[31:0] T199;
  wire[5:0] T200;
  wire T201;
  wire T202;
  wire[37:0] T203;
  wire[37:0] T204;
  wire[31:0] T205;
  wire[5:0] T206;
  wire T207;
  wire T208;
  wire[37:0] T209;
  wire[37:0] T210;
  wire[31:0] T211;
  wire[5:0] T212;
  wire T213;
  wire T214;
  wire[37:0] T215;
  wire[37:0] T216;
  wire[31:0] T217;
  wire[5:0] T218;
  wire T219;
  wire T220;
  wire[37:0] T221;
  wire[37:0] T222;
  wire[31:0] T223;
  wire[5:0] T224;
  wire T225;
  wire T226;
  wire[37:0] T227;
  wire[37:0] T228;
  wire[31:0] T229;
  wire[5:0] T230;
  wire T231;
  wire T232;
  wire[37:0] T233;
  wire[37:0] T234;
  wire[31:0] T235;
  wire[5:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  reg  nextRqstValid;
  wire T766;
  wire T242;
  wire T243;
  reg  seqInfoRegValid;
  wire T767;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire[31:0] T768;
  wire[14:0] T250;
  wire[14:0] T251;
  reg [14:0] nextRqst;
  wire[14:0] T769;
  wire[37:0] T770;
  wire[37:0] T252;
  wire[37:0] T771;
  wire[37:0] T253;
  wire[31:0] T254;
  wire[31:0] offsetAddr;
  wire[31:0] T255;
  wire[31:0] T256;
  wire[31:0] T257;
  reg [42:0] seqInfoReg;
  wire[42:0] T772;
  wire[42:0] T258;
  wire T259;
  wire[31:0] T773;
  wire[8:0] savedOffsetsVal;
  wire[8:0] T774;
  wire[31:0] T260;
  wire[31:0] T261;
  wire[31:0] T262;
  wire[31:0] T263;
  wire[31:0] T264;
  wire[31:0] T265;
  wire[31:0] T266;
  wire[31:0] spillLkup;
  wire[31:0] T267;
  wire[31:0] T268;
  wire[31:0] T775;
  wire[8:0] T579;
  wire[8:0] T580;
  wire[8:0] T581;
  wire[8:0] T582;
  wire[8:0] T583;
  reg [8:0] savedOffsets_0;
  wire[8:0] T776;
  wire[8:0] T584;
  wire[8:0] T585;
  wire T586;
  wire T587;
  wire[31:0] T588;
  wire[4:0] T589;
  wire[4:0] addrLkupIndex;
  wire[4:0] T300;
  wire[4:0] T301;
  wire[4:0] T302;
  reg [8:0] savedOffsets_1;
  wire[8:0] T777;
  wire[8:0] T590;
  wire[8:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[8:0] T595;
  reg [8:0] savedOffsets_2;
  wire[8:0] T778;
  wire[8:0] T596;
  wire[8:0] T597;
  wire T598;
  wire T599;
  reg [8:0] savedOffsets_3;
  wire[8:0] T779;
  wire[8:0] T600;
  wire[8:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire[8:0] T606;
  wire[8:0] T607;
  reg [8:0] savedOffsets_4;
  wire[8:0] T780;
  wire[8:0] T608;
  wire[8:0] T609;
  wire T610;
  wire T611;
  reg [8:0] savedOffsets_5;
  wire[8:0] T781;
  wire[8:0] T612;
  wire[8:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[8:0] T617;
  reg [8:0] savedOffsets_6;
  wire[8:0] T782;
  wire[8:0] T618;
  wire[8:0] T619;
  wire T620;
  wire T621;
  reg [8:0] savedOffsets_7;
  wire[8:0] T783;
  wire[8:0] T622;
  wire[8:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire[8:0] T629;
  wire[8:0] T630;
  wire[8:0] T631;
  reg [8:0] savedOffsets_8;
  wire[8:0] T784;
  wire[8:0] T632;
  wire[8:0] T633;
  wire T634;
  wire T635;
  reg [8:0] savedOffsets_9;
  wire[8:0] T785;
  wire[8:0] T636;
  wire[8:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[8:0] T641;
  reg [8:0] savedOffsets_10;
  wire[8:0] T786;
  wire[8:0] T642;
  wire[8:0] T643;
  wire T644;
  wire T645;
  reg [8:0] savedOffsets_11;
  wire[8:0] T787;
  wire[8:0] T646;
  wire[8:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[8:0] T652;
  wire[8:0] T653;
  reg [8:0] savedOffsets_12;
  wire[8:0] T788;
  wire[8:0] T654;
  wire[8:0] T655;
  wire T656;
  wire T657;
  reg [8:0] savedOffsets_13;
  wire[8:0] T789;
  wire[8:0] T658;
  wire[8:0] T659;
  wire T660;
  wire T661;
  wire T662;
  wire[8:0] T663;
  reg [8:0] savedOffsets_14;
  wire[8:0] T790;
  wire[8:0] T664;
  wire[8:0] T665;
  wire T666;
  wire T667;
  reg [8:0] savedOffsets_15;
  wire[8:0] T791;
  wire[8:0] T668;
  wire[8:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[8:0] T676;
  wire[8:0] T677;
  reg [8:0] savedOffsets_16;
  wire[8:0] T792;
  wire[8:0] T678;
  wire[8:0] T679;
  wire T680;
  wire T681;
  reg [8:0] savedOffsets_17;
  wire[8:0] T793;
  wire[8:0] T682;
  wire[8:0] T683;
  wire T684;
  wire T685;
  wire T686;
  wire[8:0] T687;
  reg [8:0] savedOffsets_18;
  wire[8:0] T794;
  wire[8:0] T688;
  wire[8:0] T689;
  wire T690;
  wire T691;
  reg [8:0] savedOffsets_19;
  wire[8:0] T795;
  wire[8:0] T692;
  wire[8:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T269;
  reg  epilogueAfterSpill;
  wire T796;
  wire T270;
  wire epilogueAfterSpillVal;
  wire T271;
  wire T272;
  wire spillEndVal;
  wire T273;
  wire T274;
  reg  spillEnd;
  wire T797;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire offsetUpdateVal_0;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire nextIterStartVal;
  wire T289;
  wire T290;
  reg  nextIterStart;
  wire T798;
  wire T291;
  reg  offsetUpdate_0;
  wire T799;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[31:0] T298;
  wire[4:0] T299;
  wire offsetUpdateVal_1;
  wire T303;
  wire T304;
  reg  offsetUpdate_1;
  wire T800;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire offsetUpdateVal_2;
  wire T311;
  wire T312;
  reg  offsetUpdate_2;
  wire T801;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire offsetUpdateVal_3;
  wire T317;
  wire T318;
  reg  offsetUpdate_3;
  wire T802;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire offsetUpdateVal_4;
  wire T327;
  wire T328;
  reg  offsetUpdate_4;
  wire T803;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire offsetUpdateVal_5;
  wire T333;
  wire T334;
  reg  offsetUpdate_5;
  wire T804;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire offsetUpdateVal_6;
  wire T341;
  wire T342;
  reg  offsetUpdate_6;
  wire T805;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire offsetUpdateVal_7;
  wire T347;
  wire T348;
  reg  offsetUpdate_7;
  wire T806;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire offsetUpdateVal_8;
  wire T359;
  wire T360;
  reg  offsetUpdate_8;
  wire T807;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire offsetUpdateVal_9;
  wire T365;
  wire T366;
  reg  offsetUpdate_9;
  wire T808;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire offsetUpdateVal_10;
  wire T373;
  wire T374;
  reg  offsetUpdate_10;
  wire T809;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire offsetUpdateVal_11;
  wire T379;
  wire T380;
  reg  offsetUpdate_11;
  wire T810;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire offsetUpdateVal_12;
  wire T389;
  wire T390;
  reg  offsetUpdate_12;
  wire T811;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire offsetUpdateVal_13;
  wire T395;
  wire T396;
  reg  offsetUpdate_13;
  wire T812;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire offsetUpdateVal_14;
  wire T403;
  wire T404;
  reg  offsetUpdate_14;
  wire T813;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire offsetUpdateVal_15;
  wire T409;
  wire T410;
  reg  offsetUpdate_15;
  wire T814;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire offsetUpdateVal_16;
  wire T421;
  wire T422;
  reg  offsetUpdate_16;
  wire T815;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire offsetUpdateVal_17;
  wire T427;
  wire T428;
  reg  offsetUpdate_17;
  wire T816;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire offsetUpdateVal_18;
  wire T435;
  wire T436;
  reg  offsetUpdate_18;
  wire T817;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire offsetUpdateVal_19;
  wire T441;
  wire T442;
  reg  offsetUpdate_19;
  wire T818;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire noCopyBaseAddrVal;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg  noCopyBaseAddr_0;
  wire T819;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire[31:0] T461;
  wire[4:0] T462;
  wire T463;
  wire T464;
  reg  noCopyBaseAddr_1;
  wire T820;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  reg  noCopyBaseAddr_2;
  wire T821;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  reg  noCopyBaseAddr_3;
  wire T822;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  reg  noCopyBaseAddr_4;
  wire T823;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  reg  noCopyBaseAddr_5;
  wire T824;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  reg  noCopyBaseAddr_6;
  wire T825;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  reg  noCopyBaseAddr_7;
  wire T826;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  reg  noCopyBaseAddr_8;
  wire T827;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  reg  noCopyBaseAddr_9;
  wire T828;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  reg  noCopyBaseAddr_10;
  wire T829;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  reg  noCopyBaseAddr_11;
  wire T830;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  reg  noCopyBaseAddr_12;
  wire T831;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  reg  noCopyBaseAddr_13;
  wire T832;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  reg  noCopyBaseAddr_14;
  wire T833;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  reg  noCopyBaseAddr_15;
  wire T834;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  reg  noCopyBaseAddr_16;
  wire T835;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  reg  noCopyBaseAddr_17;
  wire T836;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  reg  noCopyBaseAddr_18;
  wire T837;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  reg  noCopyBaseAddr_19;
  wire T838;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[31:0] T574;
  wire[31:0] loopOffsetLkup;
  wire[31:0] T575;
  wire[31:0] T576;
  wire[31:0] T839;
  wire T577;
  wire T578;
  wire[31:0] T840;
  wire T699;
  wire T700;
  wire[31:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire[31:0] T706;
  wire T707;
  wire T708;
  wire[31:0] baseAddrLkup;
  wire[31:0] T709;
  wire[31:0] T710;
  wire T711;
  wire T712;
  wire[5:0] nextLkupIndex;
  wire[5:0] T713;
  wire[5:0] T714;
  wire[5:0] T715;
  wire T716;
  wire lRespFifoDeq;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire[4:0] T727;
  wire T728;
  wire[4:0] T729;
  wire T730;
  wire[8:0] T731;
  wire T732;
  wire[5:0] T733;
  wire[5:0] T734;
  wire[5:0] T735;
  wire[5:0] T841;
  reg [1:0] lookupIndex;
  wire[1:0] T842;
  wire[1:0] T736;
  wire[1:0] T737;
  wire[1:0] T738;
  wire[5:0] regLookupIndex;
  wire[5:0] T739;
  wire[5:0] T740;
  wire T741;
  wire T742;
  wire[4:0] T743;
  wire T744;
  wire T745;
  wire[31:0] baseAddrMem_io_outData;
  wire[56:0] regLookupMem_io_outData;
  wire[42:0] loadSeqMem_io_outData;
  wire[31:0] loopOffsetMem_io_outData;
  wire[31:0] spillOffsetMem_io_outData;
  wire[8:0] loadSeqMemConfig_io_memAddr;
  wire[42:0] loadSeqMemConfig_io_memData;
  wire loadSeqMemConfig_io_memOutValid;
  wire loadSeqMemConfig_io_rst;
  wire[5:0] regLkupMemConfig_io_memAddr;
  wire[56:0] regLkupMemConfig_io_memData;
  wire regLkupMemConfig_io_memOutValid;
  wire[4:0] baseAddrMemConfig_io_memAddr;
  wire[31:0] baseAddrMemConfig_io_memData;
  wire baseAddrMemConfig_io_memOutValid;
  wire[4:0] loopOffsetMemConfig_io_memAddr;
  wire[31:0] loopOffsetMemConfig_io_memData;
  wire loopOffsetMemConfig_io_memOutValid;
  wire[4:0] spillOffsetMemConfig_io_memAddr;
  wire[31:0] spillOffsetMemConfig_io_memData;
  wire spillOffsetMemConfig_io_memOutValid;
  wire[37:0] lrRespFifo_io_deqData;
  wire lrRespFifo_io_enqRdy;
  wire lrRespFifo_io_deqValid;
  wire[31:0] lrReqFifo_io_deqData;
  wire lrReqFifo_io_enqRdy;
  wire lrReqFifo_io_deqValid;
  wire[37:0] fifo_io_deqData;
  wire fifo_io_enqRdy;
  wire fifo_io_deqValid;
  wire[37:0] fifo_1_io_deqData;
  wire fifo_1_io_enqRdy;
  wire fifo_1_io_deqValid;
  wire[37:0] fifo_2_io_deqData;
  wire fifo_2_io_enqRdy;
  wire fifo_2_io_deqValid;
  wire[37:0] fifo_3_io_deqData;
  wire fifo_3_io_enqRdy;
  wire fifo_3_io_deqValid;
  wire[37:0] fifo_4_io_deqData;
  wire fifo_4_io_enqRdy;
  wire fifo_4_io_deqValid;
  wire[37:0] fifo_5_io_deqData;
  wire fifo_5_io_enqRdy;
  wire fifo_5_io_deqValid;
  wire[37:0] fifo_6_io_deqData;
  wire fifo_6_io_enqRdy;
  wire fifo_6_io_deqValid;
  wire[37:0] fifo_7_io_deqData;
  wire fifo_7_io_enqRdy;
  wire fifo_7_io_deqValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lRespDest = {2{$random}};
    enqDoneReg = {1{$random}};
    lRespLkupValid = {1{$random}};
    lRespData = {1{$random}};
    nextRqstValid = {1{$random}};
    seqInfoRegValid = {1{$random}};
    nextRqst = {1{$random}};
    seqInfoReg = {2{$random}};
    savedOffsets_0 = {1{$random}};
    savedOffsets_1 = {1{$random}};
    savedOffsets_2 = {1{$random}};
    savedOffsets_3 = {1{$random}};
    savedOffsets_4 = {1{$random}};
    savedOffsets_5 = {1{$random}};
    savedOffsets_6 = {1{$random}};
    savedOffsets_7 = {1{$random}};
    savedOffsets_8 = {1{$random}};
    savedOffsets_9 = {1{$random}};
    savedOffsets_10 = {1{$random}};
    savedOffsets_11 = {1{$random}};
    savedOffsets_12 = {1{$random}};
    savedOffsets_13 = {1{$random}};
    savedOffsets_14 = {1{$random}};
    savedOffsets_15 = {1{$random}};
    savedOffsets_16 = {1{$random}};
    savedOffsets_17 = {1{$random}};
    savedOffsets_18 = {1{$random}};
    savedOffsets_19 = {1{$random}};
    epilogueAfterSpill = {1{$random}};
    spillEnd = {1{$random}};
    nextIterStart = {1{$random}};
    offsetUpdate_0 = {1{$random}};
    offsetUpdate_1 = {1{$random}};
    offsetUpdate_2 = {1{$random}};
    offsetUpdate_3 = {1{$random}};
    offsetUpdate_4 = {1{$random}};
    offsetUpdate_5 = {1{$random}};
    offsetUpdate_6 = {1{$random}};
    offsetUpdate_7 = {1{$random}};
    offsetUpdate_8 = {1{$random}};
    offsetUpdate_9 = {1{$random}};
    offsetUpdate_10 = {1{$random}};
    offsetUpdate_11 = {1{$random}};
    offsetUpdate_12 = {1{$random}};
    offsetUpdate_13 = {1{$random}};
    offsetUpdate_14 = {1{$random}};
    offsetUpdate_15 = {1{$random}};
    offsetUpdate_16 = {1{$random}};
    offsetUpdate_17 = {1{$random}};
    offsetUpdate_18 = {1{$random}};
    offsetUpdate_19 = {1{$random}};
    noCopyBaseAddr_0 = {1{$random}};
    noCopyBaseAddr_1 = {1{$random}};
    noCopyBaseAddr_2 = {1{$random}};
    noCopyBaseAddr_3 = {1{$random}};
    noCopyBaseAddr_4 = {1{$random}};
    noCopyBaseAddr_5 = {1{$random}};
    noCopyBaseAddr_6 = {1{$random}};
    noCopyBaseAddr_7 = {1{$random}};
    noCopyBaseAddr_8 = {1{$random}};
    noCopyBaseAddr_9 = {1{$random}};
    noCopyBaseAddr_10 = {1{$random}};
    noCopyBaseAddr_11 = {1{$random}};
    noCopyBaseAddr_12 = {1{$random}};
    noCopyBaseAddr_13 = {1{$random}};
    noCopyBaseAddr_14 = {1{$random}};
    noCopyBaseAddr_15 = {1{$random}};
    noCopyBaseAddr_16 = {1{$random}};
    noCopyBaseAddr_17 = {1{$random}};
    noCopyBaseAddr_18 = {1{$random}};
    noCopyBaseAddr_19 = {1{$random}};
    lookupIndex = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1 = T2 ? 1'h1 : 1'h0;
  assign T2 = enqReqWire_7 & fifo_7_io_enqRdy;
  assign enqReqWire_7 = T3;
  assign T3 = lRespLkupValid ? T4 : 1'h0;
  assign T4 = lRespDest[6'h2f:6'h2f];
  assign T746 = reset ? 57'h0 : T5;
  assign T5 = T7 ? regLookup : lRespDest;
  assign regLookup = T6;
  assign T6 = T7 ? regLookupMem_io_outData : 57'h0;
  assign T7 = lrRespFifo_io_deqValid & enqComplete;
  assign enqComplete = T8;
  assign T8 = T9;
  assign T9 = enqDoneReg == 8'hff;
  assign T747 = reset ? 8'h0 : T10;
  assign T10 = T2 ? T175 : T11;
  assign T11 = T174 ? T166 : T12;
  assign T12 = T165 ? T157 : T13;
  assign T13 = T156 ? T148 : T14;
  assign T14 = T147 ? T139 : T15;
  assign T15 = T138 ? T130 : T16;
  assign T16 = T129 ? T121 : T17;
  assign T17 = T120 ? T112 : T18;
  assign T18 = T26 | T19;
  assign T19 = T748 & T20;
  assign T20 = 8'h80 | T21;
  assign T21 = enqDoneReg ^ enqDoneReg;
  assign T748 = T22 ? 8'hff : 8'h0;
  assign T22 = T23;
  assign T23 = T24;
  assign T24 = T25 | fifo_7_io_enqRdy;
  assign T25 = ~ enqReqWire_7;
  assign T26 = T28 & T27;
  assign T27 = ~ T20;
  assign T28 = T38 | T29;
  assign T29 = T749 & T30;
  assign T30 = 8'h40 | T31;
  assign T31 = enqDoneReg ^ enqDoneReg;
  assign T749 = T32 ? 8'hff : 8'h0;
  assign T32 = T33;
  assign T33 = T34;
  assign T34 = T35 | fifo_6_io_enqRdy;
  assign T35 = ~ enqReqWire_6;
  assign enqReqWire_6 = T36;
  assign T36 = lRespLkupValid ? T37 : 1'h0;
  assign T37 = lRespDest[6'h29:6'h29];
  assign T38 = T40 & T39;
  assign T39 = ~ T30;
  assign T40 = T50 | T41;
  assign T41 = T750 & T42;
  assign T42 = 8'h20 | T43;
  assign T43 = enqDoneReg ^ enqDoneReg;
  assign T750 = T44 ? 8'hff : 8'h0;
  assign T44 = T45;
  assign T45 = T46;
  assign T46 = T47 | fifo_5_io_enqRdy;
  assign T47 = ~ enqReqWire_5;
  assign enqReqWire_5 = T48;
  assign T48 = lRespLkupValid ? T49 : 1'h0;
  assign T49 = lRespDest[6'h23:6'h23];
  assign T50 = T52 & T51;
  assign T51 = ~ T42;
  assign T52 = T62 | T53;
  assign T53 = T751 & T54;
  assign T54 = 8'h10 | T55;
  assign T55 = enqDoneReg ^ enqDoneReg;
  assign T751 = T56 ? 8'hff : 8'h0;
  assign T56 = T57;
  assign T57 = T58;
  assign T58 = T59 | fifo_4_io_enqRdy;
  assign T59 = ~ enqReqWire_4;
  assign enqReqWire_4 = T60;
  assign T60 = lRespLkupValid ? T61 : 1'h0;
  assign T61 = lRespDest[5'h1d:5'h1d];
  assign T62 = T64 & T63;
  assign T63 = ~ T54;
  assign T64 = T74 | T65;
  assign T65 = T752 & T66;
  assign T66 = 8'h8 | T67;
  assign T67 = enqDoneReg ^ enqDoneReg;
  assign T752 = T68 ? 8'hff : 8'h0;
  assign T68 = T69;
  assign T69 = T70;
  assign T70 = T71 | fifo_3_io_enqRdy;
  assign T71 = ~ enqReqWire_3;
  assign enqReqWire_3 = T72;
  assign T72 = lRespLkupValid ? T73 : 1'h0;
  assign T73 = lRespDest[5'h17:5'h17];
  assign T74 = T76 & T75;
  assign T75 = ~ T66;
  assign T76 = T86 | T77;
  assign T77 = T753 & T78;
  assign T78 = 8'h4 | T79;
  assign T79 = enqDoneReg ^ enqDoneReg;
  assign T753 = T80 ? 8'hff : 8'h0;
  assign T80 = T81;
  assign T81 = T82;
  assign T82 = T83 | fifo_2_io_enqRdy;
  assign T83 = ~ enqReqWire_2;
  assign enqReqWire_2 = T84;
  assign T84 = lRespLkupValid ? T85 : 1'h0;
  assign T85 = lRespDest[5'h11:5'h11];
  assign T86 = T88 & T87;
  assign T87 = ~ T78;
  assign T88 = T98 | T89;
  assign T89 = T754 & T90;
  assign T90 = 8'h2 | T91;
  assign T91 = enqDoneReg ^ enqDoneReg;
  assign T754 = T92 ? 8'hff : 8'h0;
  assign T92 = T93;
  assign T93 = T94;
  assign T94 = T95 | fifo_1_io_enqRdy;
  assign T95 = ~ enqReqWire_1;
  assign enqReqWire_1 = T96;
  assign T96 = lRespLkupValid ? T97 : 1'h0;
  assign T97 = lRespDest[4'hb:4'hb];
  assign T98 = T100 & T99;
  assign T99 = ~ T90;
  assign T100 = T110 | T101;
  assign T101 = T755 & T102;
  assign T102 = 8'h1 | T103;
  assign T103 = enqDoneReg ^ enqDoneReg;
  assign T755 = T104 ? 8'hff : 8'h0;
  assign T104 = T105;
  assign T105 = T106;
  assign T106 = T107 | fifo_io_enqRdy;
  assign T107 = ~ enqReqWire_0;
  assign enqReqWire_0 = T108;
  assign T108 = lRespLkupValid ? T109 : 1'h0;
  assign T109 = lRespDest[3'h5:3'h5];
  assign T110 = enqDoneReg & T111;
  assign T111 = ~ T102;
  assign T112 = T118 | T113;
  assign T113 = T756 & T114;
  assign T114 = 8'h1 | T115;
  assign T115 = enqDoneReg ^ enqDoneReg;
  assign T756 = T116 ? 8'hff : 8'h0;
  assign T116 = T117;
  assign T117 = 1'h1;
  assign T118 = T18 & T119;
  assign T119 = ~ T114;
  assign T120 = enqReqWire_0 & fifo_io_enqRdy;
  assign T121 = T127 | T122;
  assign T122 = T757 & T123;
  assign T123 = 8'h2 | T124;
  assign T124 = enqDoneReg ^ enqDoneReg;
  assign T757 = T125 ? 8'hff : 8'h0;
  assign T125 = T126;
  assign T126 = 1'h1;
  assign T127 = T17 & T128;
  assign T128 = ~ T123;
  assign T129 = enqReqWire_1 & fifo_1_io_enqRdy;
  assign T130 = T136 | T131;
  assign T131 = T758 & T132;
  assign T132 = 8'h4 | T133;
  assign T133 = enqDoneReg ^ enqDoneReg;
  assign T758 = T134 ? 8'hff : 8'h0;
  assign T134 = T135;
  assign T135 = 1'h1;
  assign T136 = T16 & T137;
  assign T137 = ~ T132;
  assign T138 = enqReqWire_2 & fifo_2_io_enqRdy;
  assign T139 = T145 | T140;
  assign T140 = T759 & T141;
  assign T141 = 8'h8 | T142;
  assign T142 = enqDoneReg ^ enqDoneReg;
  assign T759 = T143 ? 8'hff : 8'h0;
  assign T143 = T144;
  assign T144 = 1'h1;
  assign T145 = T15 & T146;
  assign T146 = ~ T141;
  assign T147 = enqReqWire_3 & fifo_3_io_enqRdy;
  assign T148 = T154 | T149;
  assign T149 = T760 & T150;
  assign T150 = 8'h10 | T151;
  assign T151 = enqDoneReg ^ enqDoneReg;
  assign T760 = T152 ? 8'hff : 8'h0;
  assign T152 = T153;
  assign T153 = 1'h1;
  assign T154 = T14 & T155;
  assign T155 = ~ T150;
  assign T156 = enqReqWire_4 & fifo_4_io_enqRdy;
  assign T157 = T163 | T158;
  assign T158 = T761 & T159;
  assign T159 = 8'h20 | T160;
  assign T160 = enqDoneReg ^ enqDoneReg;
  assign T761 = T161 ? 8'hff : 8'h0;
  assign T161 = T162;
  assign T162 = 1'h1;
  assign T163 = T13 & T164;
  assign T164 = ~ T159;
  assign T165 = enqReqWire_5 & fifo_5_io_enqRdy;
  assign T166 = T172 | T167;
  assign T167 = T762 & T168;
  assign T168 = 8'h40 | T169;
  assign T169 = enqDoneReg ^ enqDoneReg;
  assign T762 = T170 ? 8'hff : 8'h0;
  assign T170 = T171;
  assign T171 = 1'h1;
  assign T172 = T12 & T173;
  assign T173 = ~ T168;
  assign T174 = enqReqWire_6 & fifo_6_io_enqRdy;
  assign T175 = T181 | T176;
  assign T176 = T763 & T177;
  assign T177 = 8'h80 | T178;
  assign T178 = enqDoneReg ^ enqDoneReg;
  assign T763 = T179 ? 8'hff : 8'h0;
  assign T179 = T180;
  assign T180 = 1'h1;
  assign T181 = T11 & T182;
  assign T182 = ~ T177;
  assign T764 = reset ? 1'h0 : T183;
  assign T183 = T185 ? 1'h0 : T184;
  assign T184 = T7 ? 1'h1 : lRespLkupValid;
  assign T185 = T187 & T186;
  assign T186 = lrRespFifo_io_deqValid ^ 1'h1;
  assign T187 = T7 ^ 1'h1;
  assign T188 = T2 ? T189 : 38'h0;
  assign T189 = {T194, T190};
  assign T190 = lRespData[5'h1f:1'h0];
  assign T765 = reset ? 32'h0 : T191;
  assign T191 = T7 ? regLookupData : lRespData;
  assign regLookupData = T192;
  assign T192 = T7 ? T193 : 32'h0;
  assign T193 = lrRespFifo_io_deqData[5'h1f:1'h0];
  assign T194 = lRespDest[6'h36:6'h31];
  assign T195 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T196 = T174 ? 1'h1 : 1'h0;
  assign T197 = T174 ? T198 : 38'h0;
  assign T198 = {T200, T199};
  assign T199 = lRespData[5'h1f:1'h0];
  assign T200 = lRespDest[6'h2f:6'h2a];
  assign T201 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T202 = T165 ? 1'h1 : 1'h0;
  assign T203 = T165 ? T204 : 38'h0;
  assign T204 = {T206, T205};
  assign T205 = lRespData[5'h1f:1'h0];
  assign T206 = lRespDest[6'h28:6'h23];
  assign T207 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T208 = T156 ? 1'h1 : 1'h0;
  assign T209 = T156 ? T210 : 38'h0;
  assign T210 = {T212, T211};
  assign T211 = lRespData[5'h1f:1'h0];
  assign T212 = lRespDest[6'h21:5'h1c];
  assign T213 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T214 = T147 ? 1'h1 : 1'h0;
  assign T215 = T147 ? T216 : 38'h0;
  assign T216 = {T218, T217};
  assign T217 = lRespData[5'h1f:1'h0];
  assign T218 = lRespDest[5'h1a:5'h15];
  assign T219 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T220 = T138 ? 1'h1 : 1'h0;
  assign T221 = T138 ? T222 : 38'h0;
  assign T222 = {T224, T223};
  assign T223 = lRespData[5'h1f:1'h0];
  assign T224 = lRespDest[5'h13:4'he];
  assign T225 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T226 = T129 ? 1'h1 : 1'h0;
  assign T227 = T129 ? T228 : 38'h0;
  assign T228 = {T230, T229};
  assign T229 = lRespData[5'h1f:1'h0];
  assign T230 = lRespDest[4'hc:3'h7];
  assign T231 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T232 = T120 ? 1'h1 : 1'h0;
  assign T233 = T120 ? T234 : 38'h0;
  assign T234 = {T236, T235};
  assign T235 = lRespData[5'h1f:1'h0];
  assign T236 = lRespDest[3'h5:1'h0];
  assign T237 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T238 = T248 ? 1'h0 : T239;
  assign T239 = T240 ? 1'h1 : 1'h0;
  assign T240 = seqInfoRegValid & T241;
  assign T241 = nextRqstValid & lrReqFifo_io_enqRdy;
  assign T766 = reset ? 1'h0 : T242;
  assign T242 = T240 ? 1'h0 : T243;
  assign T243 = seqInfoRegValid ? 1'h1 : nextRqstValid;
  assign T767 = reset ? 1'h0 : T244;
  assign T244 = loadSeqMemConfig_io_rst ? 1'h0 : T245;
  assign T245 = seqInfoRegValid ? 1'h0 : T246;
  assign T246 = T247 ? 1'h1 : seqInfoRegValid;
  assign T247 = lrReqFifo_io_enqRdy & io_seqMemAddrValid;
  assign T248 = seqInfoRegValid & T249;
  assign T249 = T241 ^ 1'h1;
  assign T768 = {17'h0, T250};
  assign T250 = T248 ? 15'h0 : T251;
  assign T251 = T240 ? nextRqst : 15'h0;
  assign T769 = T770[4'he:1'h0];
  assign T770 = reset ? 38'h0 : T252;
  assign T252 = seqInfoRegValid ? T253 : T771;
  assign T771 = {23'h0, nextRqst};
  assign T253 = {nextLkupIndex, T254};
  assign T254 = T773 + offsetAddr;
  assign offsetAddr = T255;
  assign T255 = T259 ? 32'h0 : T256;
  assign T256 = seqInfoRegValid ? T257 : 32'h0;
  assign T257 = seqInfoReg[5'h1f:1'h0];
  assign T772 = reset ? 43'h0 : T258;
  assign T258 = T247 ? loadSeqMem_io_outData : seqInfoReg;
  assign T259 = seqInfoRegValid ^ 1'h1;
  assign T773 = {23'h0, savedOffsetsVal};
  assign savedOffsetsVal = T774;
  assign T774 = T260[4'h8:1'h0];
  assign T260 = T711 ? baseAddrLkup : T261;
  assign T261 = T707 ? T706 : T262;
  assign T262 = T702 ? T701 : T263;
  assign T263 = T699 ? T840 : T264;
  assign T264 = T577 ? T574 : T265;
  assign T265 = T269 ? T266 : 32'h0;
  assign T266 = T775 - spillLkup;
  assign spillLkup = T267;
  assign T267 = T259 ? 32'h0 : T268;
  assign T268 = seqInfoRegValid ? spillOffsetMem_io_outData : 32'h0;
  assign T775 = {23'h0, T579};
  assign T579 = T698 ? T676 : T580;
  assign T580 = T675 ? T629 : T581;
  assign T581 = T628 ? T606 : T582;
  assign T582 = T605 ? T595 : T583;
  assign T583 = T594 ? savedOffsets_1 : savedOffsets_0;
  assign T776 = reset ? 9'h0 : T584;
  assign T584 = loadSeqMemConfig_io_rst ? 9'h0 : T585;
  assign T585 = T586 ? savedOffsetsVal : savedOffsets_0;
  assign T586 = seqInfoRegValid & T587;
  assign T587 = T588[1'h0:1'h0];
  assign T588 = 1'h1 << T589;
  assign T589 = addrLkupIndex;
  assign addrLkupIndex = T300;
  assign T300 = T259 ? 5'h0 : T301;
  assign T301 = seqInfoRegValid ? T302 : 5'h0;
  assign T302 = seqInfoReg[6'h24:6'h20];
  assign T777 = reset ? 9'h0 : T590;
  assign T590 = loadSeqMemConfig_io_rst ? 9'h0 : T591;
  assign T591 = T592 ? savedOffsetsVal : savedOffsets_1;
  assign T592 = seqInfoRegValid & T593;
  assign T593 = T588[1'h1:1'h1];
  assign T594 = T589[1'h0:1'h0];
  assign T595 = T604 ? savedOffsets_3 : savedOffsets_2;
  assign T778 = reset ? 9'h0 : T596;
  assign T596 = loadSeqMemConfig_io_rst ? 9'h0 : T597;
  assign T597 = T598 ? savedOffsetsVal : savedOffsets_2;
  assign T598 = seqInfoRegValid & T599;
  assign T599 = T588[2'h2:2'h2];
  assign T779 = reset ? 9'h0 : T600;
  assign T600 = loadSeqMemConfig_io_rst ? 9'h0 : T601;
  assign T601 = T602 ? savedOffsetsVal : savedOffsets_3;
  assign T602 = seqInfoRegValid & T603;
  assign T603 = T588[2'h3:2'h3];
  assign T604 = T589[1'h0:1'h0];
  assign T605 = T589[1'h1:1'h1];
  assign T606 = T627 ? T617 : T607;
  assign T607 = T616 ? savedOffsets_5 : savedOffsets_4;
  assign T780 = reset ? 9'h0 : T608;
  assign T608 = loadSeqMemConfig_io_rst ? 9'h0 : T609;
  assign T609 = T610 ? savedOffsetsVal : savedOffsets_4;
  assign T610 = seqInfoRegValid & T611;
  assign T611 = T588[3'h4:3'h4];
  assign T781 = reset ? 9'h0 : T612;
  assign T612 = loadSeqMemConfig_io_rst ? 9'h0 : T613;
  assign T613 = T614 ? savedOffsetsVal : savedOffsets_5;
  assign T614 = seqInfoRegValid & T615;
  assign T615 = T588[3'h5:3'h5];
  assign T616 = T589[1'h0:1'h0];
  assign T617 = T626 ? savedOffsets_7 : savedOffsets_6;
  assign T782 = reset ? 9'h0 : T618;
  assign T618 = loadSeqMemConfig_io_rst ? 9'h0 : T619;
  assign T619 = T620 ? savedOffsetsVal : savedOffsets_6;
  assign T620 = seqInfoRegValid & T621;
  assign T621 = T588[3'h6:3'h6];
  assign T783 = reset ? 9'h0 : T622;
  assign T622 = loadSeqMemConfig_io_rst ? 9'h0 : T623;
  assign T623 = T624 ? savedOffsetsVal : savedOffsets_7;
  assign T624 = seqInfoRegValid & T625;
  assign T625 = T588[3'h7:3'h7];
  assign T626 = T589[1'h0:1'h0];
  assign T627 = T589[1'h1:1'h1];
  assign T628 = T589[2'h2:2'h2];
  assign T629 = T674 ? T652 : T630;
  assign T630 = T651 ? T641 : T631;
  assign T631 = T640 ? savedOffsets_9 : savedOffsets_8;
  assign T784 = reset ? 9'h0 : T632;
  assign T632 = loadSeqMemConfig_io_rst ? 9'h0 : T633;
  assign T633 = T634 ? savedOffsetsVal : savedOffsets_8;
  assign T634 = seqInfoRegValid & T635;
  assign T635 = T588[4'h8:4'h8];
  assign T785 = reset ? 9'h0 : T636;
  assign T636 = loadSeqMemConfig_io_rst ? 9'h0 : T637;
  assign T637 = T638 ? savedOffsetsVal : savedOffsets_9;
  assign T638 = seqInfoRegValid & T639;
  assign T639 = T588[4'h9:4'h9];
  assign T640 = T589[1'h0:1'h0];
  assign T641 = T650 ? savedOffsets_11 : savedOffsets_10;
  assign T786 = reset ? 9'h0 : T642;
  assign T642 = loadSeqMemConfig_io_rst ? 9'h0 : T643;
  assign T643 = T644 ? savedOffsetsVal : savedOffsets_10;
  assign T644 = seqInfoRegValid & T645;
  assign T645 = T588[4'ha:4'ha];
  assign T787 = reset ? 9'h0 : T646;
  assign T646 = loadSeqMemConfig_io_rst ? 9'h0 : T647;
  assign T647 = T648 ? savedOffsetsVal : savedOffsets_11;
  assign T648 = seqInfoRegValid & T649;
  assign T649 = T588[4'hb:4'hb];
  assign T650 = T589[1'h0:1'h0];
  assign T651 = T589[1'h1:1'h1];
  assign T652 = T673 ? T663 : T653;
  assign T653 = T662 ? savedOffsets_13 : savedOffsets_12;
  assign T788 = reset ? 9'h0 : T654;
  assign T654 = loadSeqMemConfig_io_rst ? 9'h0 : T655;
  assign T655 = T656 ? savedOffsetsVal : savedOffsets_12;
  assign T656 = seqInfoRegValid & T657;
  assign T657 = T588[4'hc:4'hc];
  assign T789 = reset ? 9'h0 : T658;
  assign T658 = loadSeqMemConfig_io_rst ? 9'h0 : T659;
  assign T659 = T660 ? savedOffsetsVal : savedOffsets_13;
  assign T660 = seqInfoRegValid & T661;
  assign T661 = T588[4'hd:4'hd];
  assign T662 = T589[1'h0:1'h0];
  assign T663 = T672 ? savedOffsets_15 : savedOffsets_14;
  assign T790 = reset ? 9'h0 : T664;
  assign T664 = loadSeqMemConfig_io_rst ? 9'h0 : T665;
  assign T665 = T666 ? savedOffsetsVal : savedOffsets_14;
  assign T666 = seqInfoRegValid & T667;
  assign T667 = T588[4'he:4'he];
  assign T791 = reset ? 9'h0 : T668;
  assign T668 = loadSeqMemConfig_io_rst ? 9'h0 : T669;
  assign T669 = T670 ? savedOffsetsVal : savedOffsets_15;
  assign T670 = seqInfoRegValid & T671;
  assign T671 = T588[4'hf:4'hf];
  assign T672 = T589[1'h0:1'h0];
  assign T673 = T589[1'h1:1'h1];
  assign T674 = T589[2'h2:2'h2];
  assign T675 = T589[2'h3:2'h3];
  assign T676 = T697 ? T687 : T677;
  assign T677 = T686 ? savedOffsets_17 : savedOffsets_16;
  assign T792 = reset ? 9'h0 : T678;
  assign T678 = loadSeqMemConfig_io_rst ? 9'h0 : T679;
  assign T679 = T680 ? savedOffsetsVal : savedOffsets_16;
  assign T680 = seqInfoRegValid & T681;
  assign T681 = T588[5'h10:5'h10];
  assign T793 = reset ? 9'h0 : T682;
  assign T682 = loadSeqMemConfig_io_rst ? 9'h0 : T683;
  assign T683 = T684 ? savedOffsetsVal : savedOffsets_17;
  assign T684 = seqInfoRegValid & T685;
  assign T685 = T588[5'h11:5'h11];
  assign T686 = T589[1'h0:1'h0];
  assign T687 = T696 ? savedOffsets_19 : savedOffsets_18;
  assign T794 = reset ? 9'h0 : T688;
  assign T688 = loadSeqMemConfig_io_rst ? 9'h0 : T689;
  assign T689 = T690 ? savedOffsetsVal : savedOffsets_18;
  assign T690 = seqInfoRegValid & T691;
  assign T691 = T588[5'h12:5'h12];
  assign T795 = reset ? 9'h0 : T692;
  assign T692 = loadSeqMemConfig_io_rst ? 9'h0 : T693;
  assign T693 = T694 ? savedOffsetsVal : savedOffsets_19;
  assign T694 = seqInfoRegValid & T695;
  assign T695 = T588[5'h13:5'h13];
  assign T696 = T589[1'h0:1'h0];
  assign T697 = T589[1'h1:1'h1];
  assign T698 = T589[3'h4:3'h4];
  assign T269 = T279 & epilogueAfterSpill;
  assign T796 = reset ? 1'h0 : T270;
  assign T270 = seqInfoRegValid ? epilogueAfterSpillVal : epilogueAfterSpill;
  assign epilogueAfterSpillVal = T271;
  assign T271 = T277 ? epilogueAfterSpill : T272;
  assign T272 = seqInfoRegValid & spillEndVal;
  assign spillEndVal = T273;
  assign T273 = T259 ? 1'h0 : T274;
  assign T274 = seqInfoRegValid ? spillEnd : 1'h0;
  assign T797 = reset ? 1'h0 : T275;
  assign T275 = loadSeqMemConfig_io_rst ? 1'h0 : T276;
  assign T276 = T247 ? io_spillEnd : spillEnd;
  assign T277 = seqInfoRegValid & T278;
  assign T278 = spillEndVal ^ 1'h1;
  assign T279 = T450 & T280;
  assign T280 = T449 ? T419 : T281;
  assign T281 = T418 ? T356 : T282;
  assign T282 = T355 ? T325 : T283;
  assign T283 = T324 ? T310 : T284;
  assign T284 = T309 ? offsetUpdateVal_1 : offsetUpdateVal_0;
  assign offsetUpdateVal_0 = T285;
  assign T285 = T296 ? 1'h0 : T286;
  assign T286 = T294 ? offsetUpdate_0 : T287;
  assign T287 = seqInfoRegValid & T288;
  assign T288 = spillEndVal | nextIterStartVal;
  assign nextIterStartVal = T289;
  assign T289 = T259 ? 1'h0 : T290;
  assign T290 = seqInfoRegValid ? nextIterStart : 1'h0;
  assign T798 = reset ? 1'h0 : T291;
  assign T291 = T247 ? io_nextIterStart : nextIterStart;
  assign T799 = reset ? 1'h0 : T292;
  assign T292 = loadSeqMemConfig_io_rst ? 1'h0 : T293;
  assign T293 = seqInfoRegValid ? offsetUpdateVal_0 : offsetUpdate_0;
  assign T294 = seqInfoRegValid & T295;
  assign T295 = T288 ^ 1'h1;
  assign T296 = seqInfoRegValid & T297;
  assign T297 = T298[1'h0:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = addrLkupIndex;
  assign offsetUpdateVal_1 = T303;
  assign T303 = T307 ? 1'h0 : T304;
  assign T304 = T294 ? offsetUpdate_1 : T287;
  assign T800 = reset ? 1'h0 : T305;
  assign T305 = loadSeqMemConfig_io_rst ? 1'h0 : T306;
  assign T306 = seqInfoRegValid ? offsetUpdateVal_1 : offsetUpdate_1;
  assign T307 = seqInfoRegValid & T308;
  assign T308 = T298[1'h1:1'h1];
  assign T309 = T299[1'h0:1'h0];
  assign T310 = T323 ? offsetUpdateVal_3 : offsetUpdateVal_2;
  assign offsetUpdateVal_2 = T311;
  assign T311 = T315 ? 1'h0 : T312;
  assign T312 = T294 ? offsetUpdate_2 : T287;
  assign T801 = reset ? 1'h0 : T313;
  assign T313 = loadSeqMemConfig_io_rst ? 1'h0 : T314;
  assign T314 = seqInfoRegValid ? offsetUpdateVal_2 : offsetUpdate_2;
  assign T315 = seqInfoRegValid & T316;
  assign T316 = T298[2'h2:2'h2];
  assign offsetUpdateVal_3 = T317;
  assign T317 = T321 ? 1'h0 : T318;
  assign T318 = T294 ? offsetUpdate_3 : T287;
  assign T802 = reset ? 1'h0 : T319;
  assign T319 = loadSeqMemConfig_io_rst ? 1'h0 : T320;
  assign T320 = seqInfoRegValid ? offsetUpdateVal_3 : offsetUpdate_3;
  assign T321 = seqInfoRegValid & T322;
  assign T322 = T298[2'h3:2'h3];
  assign T323 = T299[1'h0:1'h0];
  assign T324 = T299[1'h1:1'h1];
  assign T325 = T354 ? T340 : T326;
  assign T326 = T339 ? offsetUpdateVal_5 : offsetUpdateVal_4;
  assign offsetUpdateVal_4 = T327;
  assign T327 = T331 ? 1'h0 : T328;
  assign T328 = T294 ? offsetUpdate_4 : T287;
  assign T803 = reset ? 1'h0 : T329;
  assign T329 = loadSeqMemConfig_io_rst ? 1'h0 : T330;
  assign T330 = seqInfoRegValid ? offsetUpdateVal_4 : offsetUpdate_4;
  assign T331 = seqInfoRegValid & T332;
  assign T332 = T298[3'h4:3'h4];
  assign offsetUpdateVal_5 = T333;
  assign T333 = T337 ? 1'h0 : T334;
  assign T334 = T294 ? offsetUpdate_5 : T287;
  assign T804 = reset ? 1'h0 : T335;
  assign T335 = loadSeqMemConfig_io_rst ? 1'h0 : T336;
  assign T336 = seqInfoRegValid ? offsetUpdateVal_5 : offsetUpdate_5;
  assign T337 = seqInfoRegValid & T338;
  assign T338 = T298[3'h5:3'h5];
  assign T339 = T299[1'h0:1'h0];
  assign T340 = T353 ? offsetUpdateVal_7 : offsetUpdateVal_6;
  assign offsetUpdateVal_6 = T341;
  assign T341 = T345 ? 1'h0 : T342;
  assign T342 = T294 ? offsetUpdate_6 : T287;
  assign T805 = reset ? 1'h0 : T343;
  assign T343 = loadSeqMemConfig_io_rst ? 1'h0 : T344;
  assign T344 = seqInfoRegValid ? offsetUpdateVal_6 : offsetUpdate_6;
  assign T345 = seqInfoRegValid & T346;
  assign T346 = T298[3'h6:3'h6];
  assign offsetUpdateVal_7 = T347;
  assign T347 = T351 ? 1'h0 : T348;
  assign T348 = T294 ? offsetUpdate_7 : T287;
  assign T806 = reset ? 1'h0 : T349;
  assign T349 = loadSeqMemConfig_io_rst ? 1'h0 : T350;
  assign T350 = seqInfoRegValid ? offsetUpdateVal_7 : offsetUpdate_7;
  assign T351 = seqInfoRegValid & T352;
  assign T352 = T298[3'h7:3'h7];
  assign T353 = T299[1'h0:1'h0];
  assign T354 = T299[1'h1:1'h1];
  assign T355 = T299[2'h2:2'h2];
  assign T356 = T417 ? T387 : T357;
  assign T357 = T386 ? T372 : T358;
  assign T358 = T371 ? offsetUpdateVal_9 : offsetUpdateVal_8;
  assign offsetUpdateVal_8 = T359;
  assign T359 = T363 ? 1'h0 : T360;
  assign T360 = T294 ? offsetUpdate_8 : T287;
  assign T807 = reset ? 1'h0 : T361;
  assign T361 = loadSeqMemConfig_io_rst ? 1'h0 : T362;
  assign T362 = seqInfoRegValid ? offsetUpdateVal_8 : offsetUpdate_8;
  assign T363 = seqInfoRegValid & T364;
  assign T364 = T298[4'h8:4'h8];
  assign offsetUpdateVal_9 = T365;
  assign T365 = T369 ? 1'h0 : T366;
  assign T366 = T294 ? offsetUpdate_9 : T287;
  assign T808 = reset ? 1'h0 : T367;
  assign T367 = loadSeqMemConfig_io_rst ? 1'h0 : T368;
  assign T368 = seqInfoRegValid ? offsetUpdateVal_9 : offsetUpdate_9;
  assign T369 = seqInfoRegValid & T370;
  assign T370 = T298[4'h9:4'h9];
  assign T371 = T299[1'h0:1'h0];
  assign T372 = T385 ? offsetUpdateVal_11 : offsetUpdateVal_10;
  assign offsetUpdateVal_10 = T373;
  assign T373 = T377 ? 1'h0 : T374;
  assign T374 = T294 ? offsetUpdate_10 : T287;
  assign T809 = reset ? 1'h0 : T375;
  assign T375 = loadSeqMemConfig_io_rst ? 1'h0 : T376;
  assign T376 = seqInfoRegValid ? offsetUpdateVal_10 : offsetUpdate_10;
  assign T377 = seqInfoRegValid & T378;
  assign T378 = T298[4'ha:4'ha];
  assign offsetUpdateVal_11 = T379;
  assign T379 = T383 ? 1'h0 : T380;
  assign T380 = T294 ? offsetUpdate_11 : T287;
  assign T810 = reset ? 1'h0 : T381;
  assign T381 = loadSeqMemConfig_io_rst ? 1'h0 : T382;
  assign T382 = seqInfoRegValid ? offsetUpdateVal_11 : offsetUpdate_11;
  assign T383 = seqInfoRegValid & T384;
  assign T384 = T298[4'hb:4'hb];
  assign T385 = T299[1'h0:1'h0];
  assign T386 = T299[1'h1:1'h1];
  assign T387 = T416 ? T402 : T388;
  assign T388 = T401 ? offsetUpdateVal_13 : offsetUpdateVal_12;
  assign offsetUpdateVal_12 = T389;
  assign T389 = T393 ? 1'h0 : T390;
  assign T390 = T294 ? offsetUpdate_12 : T287;
  assign T811 = reset ? 1'h0 : T391;
  assign T391 = loadSeqMemConfig_io_rst ? 1'h0 : T392;
  assign T392 = seqInfoRegValid ? offsetUpdateVal_12 : offsetUpdate_12;
  assign T393 = seqInfoRegValid & T394;
  assign T394 = T298[4'hc:4'hc];
  assign offsetUpdateVal_13 = T395;
  assign T395 = T399 ? 1'h0 : T396;
  assign T396 = T294 ? offsetUpdate_13 : T287;
  assign T812 = reset ? 1'h0 : T397;
  assign T397 = loadSeqMemConfig_io_rst ? 1'h0 : T398;
  assign T398 = seqInfoRegValid ? offsetUpdateVal_13 : offsetUpdate_13;
  assign T399 = seqInfoRegValid & T400;
  assign T400 = T298[4'hd:4'hd];
  assign T401 = T299[1'h0:1'h0];
  assign T402 = T415 ? offsetUpdateVal_15 : offsetUpdateVal_14;
  assign offsetUpdateVal_14 = T403;
  assign T403 = T407 ? 1'h0 : T404;
  assign T404 = T294 ? offsetUpdate_14 : T287;
  assign T813 = reset ? 1'h0 : T405;
  assign T405 = loadSeqMemConfig_io_rst ? 1'h0 : T406;
  assign T406 = seqInfoRegValid ? offsetUpdateVal_14 : offsetUpdate_14;
  assign T407 = seqInfoRegValid & T408;
  assign T408 = T298[4'he:4'he];
  assign offsetUpdateVal_15 = T409;
  assign T409 = T413 ? 1'h0 : T410;
  assign T410 = T294 ? offsetUpdate_15 : T287;
  assign T814 = reset ? 1'h0 : T411;
  assign T411 = loadSeqMemConfig_io_rst ? 1'h0 : T412;
  assign T412 = seqInfoRegValid ? offsetUpdateVal_15 : offsetUpdate_15;
  assign T413 = seqInfoRegValid & T414;
  assign T414 = T298[4'hf:4'hf];
  assign T415 = T299[1'h0:1'h0];
  assign T416 = T299[1'h1:1'h1];
  assign T417 = T299[2'h2:2'h2];
  assign T418 = T299[2'h3:2'h3];
  assign T419 = T448 ? T434 : T420;
  assign T420 = T433 ? offsetUpdateVal_17 : offsetUpdateVal_16;
  assign offsetUpdateVal_16 = T421;
  assign T421 = T425 ? 1'h0 : T422;
  assign T422 = T294 ? offsetUpdate_16 : T287;
  assign T815 = reset ? 1'h0 : T423;
  assign T423 = loadSeqMemConfig_io_rst ? 1'h0 : T424;
  assign T424 = seqInfoRegValid ? offsetUpdateVal_16 : offsetUpdate_16;
  assign T425 = seqInfoRegValid & T426;
  assign T426 = T298[5'h10:5'h10];
  assign offsetUpdateVal_17 = T427;
  assign T427 = T431 ? 1'h0 : T428;
  assign T428 = T294 ? offsetUpdate_17 : T287;
  assign T816 = reset ? 1'h0 : T429;
  assign T429 = loadSeqMemConfig_io_rst ? 1'h0 : T430;
  assign T430 = seqInfoRegValid ? offsetUpdateVal_17 : offsetUpdate_17;
  assign T431 = seqInfoRegValid & T432;
  assign T432 = T298[5'h11:5'h11];
  assign T433 = T299[1'h0:1'h0];
  assign T434 = T447 ? offsetUpdateVal_19 : offsetUpdateVal_18;
  assign offsetUpdateVal_18 = T435;
  assign T435 = T439 ? 1'h0 : T436;
  assign T436 = T294 ? offsetUpdate_18 : T287;
  assign T817 = reset ? 1'h0 : T437;
  assign T437 = loadSeqMemConfig_io_rst ? 1'h0 : T438;
  assign T438 = seqInfoRegValid ? offsetUpdateVal_18 : offsetUpdate_18;
  assign T439 = seqInfoRegValid & T440;
  assign T440 = T298[5'h12:5'h12];
  assign offsetUpdateVal_19 = T441;
  assign T441 = T445 ? 1'h0 : T442;
  assign T442 = T294 ? offsetUpdate_19 : T287;
  assign T818 = reset ? 1'h0 : T443;
  assign T443 = loadSeqMemConfig_io_rst ? 1'h0 : T444;
  assign T444 = seqInfoRegValid ? offsetUpdateVal_19 : offsetUpdate_19;
  assign T445 = seqInfoRegValid & T446;
  assign T446 = T298[5'h13:5'h13];
  assign T447 = T299[1'h0:1'h0];
  assign T448 = T299[1'h1:1'h1];
  assign T449 = T299[3'h4:3'h4];
  assign T450 = seqInfoRegValid & noCopyBaseAddrVal;
  assign noCopyBaseAddrVal = T451;
  assign T451 = seqInfoRegValid ? T452 : 1'h0;
  assign T452 = T573 ? T551 : T453;
  assign T453 = T550 ? T504 : T454;
  assign T454 = T503 ? T481 : T455;
  assign T455 = T480 ? T470 : T456;
  assign T456 = T469 ? noCopyBaseAddr_1 : noCopyBaseAddr_0;
  assign T819 = reset ? 1'h0 : T457;
  assign T457 = loadSeqMemConfig_io_rst ? 1'h0 : T458;
  assign T458 = T459 ? 1'h1 : noCopyBaseAddr_0;
  assign T459 = T463 & T460;
  assign T460 = T461[1'h0:1'h0];
  assign T461 = 1'h1 << T462;
  assign T462 = addrLkupIndex;
  assign T463 = seqInfoRegValid & T464;
  assign T464 = noCopyBaseAddrVal ^ 1'h1;
  assign T820 = reset ? 1'h0 : T465;
  assign T465 = loadSeqMemConfig_io_rst ? 1'h0 : T466;
  assign T466 = T467 ? 1'h1 : noCopyBaseAddr_1;
  assign T467 = T463 & T468;
  assign T468 = T461[1'h1:1'h1];
  assign T469 = T462[1'h0:1'h0];
  assign T470 = T479 ? noCopyBaseAddr_3 : noCopyBaseAddr_2;
  assign T821 = reset ? 1'h0 : T471;
  assign T471 = loadSeqMemConfig_io_rst ? 1'h0 : T472;
  assign T472 = T473 ? 1'h1 : noCopyBaseAddr_2;
  assign T473 = T463 & T474;
  assign T474 = T461[2'h2:2'h2];
  assign T822 = reset ? 1'h0 : T475;
  assign T475 = loadSeqMemConfig_io_rst ? 1'h0 : T476;
  assign T476 = T477 ? 1'h1 : noCopyBaseAddr_3;
  assign T477 = T463 & T478;
  assign T478 = T461[2'h3:2'h3];
  assign T479 = T462[1'h0:1'h0];
  assign T480 = T462[1'h1:1'h1];
  assign T481 = T502 ? T492 : T482;
  assign T482 = T491 ? noCopyBaseAddr_5 : noCopyBaseAddr_4;
  assign T823 = reset ? 1'h0 : T483;
  assign T483 = loadSeqMemConfig_io_rst ? 1'h0 : T484;
  assign T484 = T485 ? 1'h1 : noCopyBaseAddr_4;
  assign T485 = T463 & T486;
  assign T486 = T461[3'h4:3'h4];
  assign T824 = reset ? 1'h0 : T487;
  assign T487 = loadSeqMemConfig_io_rst ? 1'h0 : T488;
  assign T488 = T489 ? 1'h1 : noCopyBaseAddr_5;
  assign T489 = T463 & T490;
  assign T490 = T461[3'h5:3'h5];
  assign T491 = T462[1'h0:1'h0];
  assign T492 = T501 ? noCopyBaseAddr_7 : noCopyBaseAddr_6;
  assign T825 = reset ? 1'h0 : T493;
  assign T493 = loadSeqMemConfig_io_rst ? 1'h0 : T494;
  assign T494 = T495 ? 1'h1 : noCopyBaseAddr_6;
  assign T495 = T463 & T496;
  assign T496 = T461[3'h6:3'h6];
  assign T826 = reset ? 1'h0 : T497;
  assign T497 = loadSeqMemConfig_io_rst ? 1'h0 : T498;
  assign T498 = T499 ? 1'h1 : noCopyBaseAddr_7;
  assign T499 = T463 & T500;
  assign T500 = T461[3'h7:3'h7];
  assign T501 = T462[1'h0:1'h0];
  assign T502 = T462[1'h1:1'h1];
  assign T503 = T462[2'h2:2'h2];
  assign T504 = T549 ? T527 : T505;
  assign T505 = T526 ? T516 : T506;
  assign T506 = T515 ? noCopyBaseAddr_9 : noCopyBaseAddr_8;
  assign T827 = reset ? 1'h0 : T507;
  assign T507 = loadSeqMemConfig_io_rst ? 1'h0 : T508;
  assign T508 = T509 ? 1'h1 : noCopyBaseAddr_8;
  assign T509 = T463 & T510;
  assign T510 = T461[4'h8:4'h8];
  assign T828 = reset ? 1'h0 : T511;
  assign T511 = loadSeqMemConfig_io_rst ? 1'h0 : T512;
  assign T512 = T513 ? 1'h1 : noCopyBaseAddr_9;
  assign T513 = T463 & T514;
  assign T514 = T461[4'h9:4'h9];
  assign T515 = T462[1'h0:1'h0];
  assign T516 = T525 ? noCopyBaseAddr_11 : noCopyBaseAddr_10;
  assign T829 = reset ? 1'h0 : T517;
  assign T517 = loadSeqMemConfig_io_rst ? 1'h0 : T518;
  assign T518 = T519 ? 1'h1 : noCopyBaseAddr_10;
  assign T519 = T463 & T520;
  assign T520 = T461[4'ha:4'ha];
  assign T830 = reset ? 1'h0 : T521;
  assign T521 = loadSeqMemConfig_io_rst ? 1'h0 : T522;
  assign T522 = T523 ? 1'h1 : noCopyBaseAddr_11;
  assign T523 = T463 & T524;
  assign T524 = T461[4'hb:4'hb];
  assign T525 = T462[1'h0:1'h0];
  assign T526 = T462[1'h1:1'h1];
  assign T527 = T548 ? T538 : T528;
  assign T528 = T537 ? noCopyBaseAddr_13 : noCopyBaseAddr_12;
  assign T831 = reset ? 1'h0 : T529;
  assign T529 = loadSeqMemConfig_io_rst ? 1'h0 : T530;
  assign T530 = T531 ? 1'h1 : noCopyBaseAddr_12;
  assign T531 = T463 & T532;
  assign T532 = T461[4'hc:4'hc];
  assign T832 = reset ? 1'h0 : T533;
  assign T533 = loadSeqMemConfig_io_rst ? 1'h0 : T534;
  assign T534 = T535 ? 1'h1 : noCopyBaseAddr_13;
  assign T535 = T463 & T536;
  assign T536 = T461[4'hd:4'hd];
  assign T537 = T462[1'h0:1'h0];
  assign T538 = T547 ? noCopyBaseAddr_15 : noCopyBaseAddr_14;
  assign T833 = reset ? 1'h0 : T539;
  assign T539 = loadSeqMemConfig_io_rst ? 1'h0 : T540;
  assign T540 = T541 ? 1'h1 : noCopyBaseAddr_14;
  assign T541 = T463 & T542;
  assign T542 = T461[4'he:4'he];
  assign T834 = reset ? 1'h0 : T543;
  assign T543 = loadSeqMemConfig_io_rst ? 1'h0 : T544;
  assign T544 = T545 ? 1'h1 : noCopyBaseAddr_15;
  assign T545 = T463 & T546;
  assign T546 = T461[4'hf:4'hf];
  assign T547 = T462[1'h0:1'h0];
  assign T548 = T462[1'h1:1'h1];
  assign T549 = T462[2'h2:2'h2];
  assign T550 = T462[2'h3:2'h3];
  assign T551 = T572 ? T562 : T552;
  assign T552 = T561 ? noCopyBaseAddr_17 : noCopyBaseAddr_16;
  assign T835 = reset ? 1'h0 : T553;
  assign T553 = loadSeqMemConfig_io_rst ? 1'h0 : T554;
  assign T554 = T555 ? 1'h1 : noCopyBaseAddr_16;
  assign T555 = T463 & T556;
  assign T556 = T461[5'h10:5'h10];
  assign T836 = reset ? 1'h0 : T557;
  assign T557 = loadSeqMemConfig_io_rst ? 1'h0 : T558;
  assign T558 = T559 ? 1'h1 : noCopyBaseAddr_17;
  assign T559 = T463 & T560;
  assign T560 = T461[5'h11:5'h11];
  assign T561 = T462[1'h0:1'h0];
  assign T562 = T571 ? noCopyBaseAddr_19 : noCopyBaseAddr_18;
  assign T837 = reset ? 1'h0 : T563;
  assign T563 = loadSeqMemConfig_io_rst ? 1'h0 : T564;
  assign T564 = T565 ? 1'h1 : noCopyBaseAddr_18;
  assign T565 = T463 & T566;
  assign T566 = T461[5'h12:5'h12];
  assign T838 = reset ? 1'h0 : T567;
  assign T567 = loadSeqMemConfig_io_rst ? 1'h0 : T568;
  assign T568 = T569 ? 1'h1 : noCopyBaseAddr_19;
  assign T569 = T463 & T570;
  assign T570 = T461[5'h13:5'h13];
  assign T571 = T462[1'h0:1'h0];
  assign T572 = T462[1'h1:1'h1];
  assign T573 = T462[3'h4:3'h4];
  assign T574 = T839 + loopOffsetLkup;
  assign loopOffsetLkup = T575;
  assign T575 = T259 ? 32'h0 : T576;
  assign T576 = seqInfoRegValid ? loopOffsetMem_io_outData : 32'h0;
  assign T839 = {23'h0, T579};
  assign T577 = T279 & T578;
  assign T578 = epilogueAfterSpill ^ 1'h1;
  assign T840 = {23'h0, T579};
  assign T699 = T450 & T700;
  assign T700 = T280 ^ 1'h1;
  assign T701 = baseAddrLkup - spillLkup;
  assign T702 = T703 & epilogueAfterSpill;
  assign T703 = T704 & T280;
  assign T704 = seqInfoRegValid & T705;
  assign T705 = noCopyBaseAddrVal ^ 1'h1;
  assign T706 = baseAddrLkup + loopOffsetLkup;
  assign T707 = T703 & T708;
  assign T708 = epilogueAfterSpill ^ 1'h1;
  assign baseAddrLkup = T709;
  assign T709 = T259 ? 32'h0 : T710;
  assign T710 = seqInfoRegValid ? baseAddrMem_io_outData : 32'h0;
  assign T711 = T704 & T712;
  assign T712 = T280 ^ 1'h1;
  assign nextLkupIndex = T713;
  assign T713 = T259 ? 6'h0 : T714;
  assign T714 = seqInfoRegValid ? T715 : 6'h0;
  assign T715 = seqInfoReg[6'h2a:6'h25];
  assign T716 = loadSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign lRespFifoDeq = T717;
  assign T717 = T725 ? 1'h0 : T718;
  assign T718 = T185 ? 1'h0 : T719;
  assign T719 = T723 ? 1'h0 : T720;
  assign T720 = T7 & T721;
  assign T721 = T722 == 1'h1;
  assign T722 = regLookup[6'h38:6'h38];
  assign T723 = T7 & T724;
  assign T724 = T721 ^ 1'h1;
  assign T725 = T726 ^ 1'h1;
  assign T726 = T7 | T186;
  assign T727 = seqInfoRegValid ? addrLkupIndex : 5'h0;
  assign T728 = seqInfoRegValid ? 1'h1 : 1'h1;
  assign T729 = seqInfoRegValid ? addrLkupIndex : 5'h0;
  assign T730 = seqInfoRegValid ? 1'h1 : 1'h1;
  assign T731 = T247 ? io_seqMemAddr : 9'h0;
  assign T732 = T247 ? io_seqMemAddrValid : 1'h0;
  assign T733 = T185 ? 6'h0 : T734;
  assign T734 = T7 ? T735 : 6'h0;
  assign T735 = regLookupIndex + T841;
  assign T841 = {4'h0, lookupIndex};
  assign T842 = reset ? 2'h0 : T736;
  assign T736 = T723 ? T738 : T737;
  assign T737 = T720 ? 2'h0 : lookupIndex;
  assign T738 = lookupIndex + 2'h1;
  assign regLookupIndex = T739;
  assign T739 = T7 ? T740 : 6'h0;
  assign T740 = lrRespFifo_io_deqData[6'h25:6'h20];
  assign T741 = T185 ? 1'h0 : T742;
  assign T742 = T7 ? 1'h1 : 1'h0;
  assign T743 = seqInfoRegValid ? addrLkupIndex : 5'h0;
  assign T744 = seqInfoRegValid ? 1'h1 : 1'h0;
  assign io_seqProceed = T745;
  assign T745 = T247 ? 1'h1 : 1'h0;
  assign io_loadRespRdy = lrRespFifo_io_enqRdy;
  assign io_loadRqstValid = lrReqFifo_io_deqValid;
  assign io_loadRqst = lrReqFifo_io_deqData;
  assign io_memBankValid_0 = fifo_io_deqValid;
  assign io_memBankValid_1 = fifo_1_io_deqValid;
  assign io_memBankValid_2 = fifo_2_io_deqValid;
  assign io_memBankValid_3 = fifo_3_io_deqValid;
  assign io_memBankValid_4 = fifo_4_io_deqValid;
  assign io_memBankValid_5 = fifo_5_io_deqValid;
  assign io_memBankValid_6 = fifo_6_io_deqValid;
  assign io_memBankValid_7 = fifo_7_io_deqValid;
  assign io_memBankEnq_0 = fifo_io_deqData;
  assign io_memBankEnq_1 = fifo_1_io_deqData;
  assign io_memBankEnq_2 = fifo_2_io_deqData;
  assign io_memBankEnq_3 = fifo_3_io_deqData;
  assign io_memBankEnq_4 = fifo_4_io_deqData;
  assign io_memBankEnq_5 = fifo_5_io_deqData;
  assign io_memBankEnq_6 = fifo_6_io_deqData;
  assign io_memBankEnq_7 = fifo_7_io_deqData;
  customReg_1 baseAddrMem(.clk(clk),
       .io_inData( baseAddrMemConfig_io_memData ),
       .io_outData( baseAddrMem_io_outData ),
       .io_readEn( T744 ),
       .io_writeEn( baseAddrMemConfig_io_memOutValid ),
       .io_readAddr( T743 ),
       .io_writeAddr( baseAddrMemConfig_io_memAddr )
  );
  customReg_2 regLookupMem(.clk(clk),
       .io_inData( regLkupMemConfig_io_memData ),
       .io_outData( regLookupMem_io_outData ),
       .io_readEn( T741 ),
       .io_writeEn( regLkupMemConfig_io_memOutValid ),
       .io_readAddr( T733 ),
       .io_writeAddr( regLkupMemConfig_io_memAddr )
  );
  customReg_3 loadSeqMem(.clk(clk),
       .io_inData( loadSeqMemConfig_io_memData ),
       .io_outData( loadSeqMem_io_outData ),
       .io_readEn( T732 ),
       .io_writeEn( loadSeqMemConfig_io_memOutValid ),
       .io_readAddr( T731 ),
       .io_writeAddr( loadSeqMemConfig_io_memAddr )
  );
  customReg_1 loopOffsetMem(.clk(clk),
       .io_inData( loopOffsetMemConfig_io_memData ),
       .io_outData( loopOffsetMem_io_outData ),
       .io_readEn( T730 ),
       .io_writeEn( loopOffsetMemConfig_io_memOutValid ),
       .io_readAddr( T729 ),
       .io_writeAddr( loopOffsetMemConfig_io_memAddr )
  );
  customReg_1 spillOffsetMem(.clk(clk),
       .io_inData( spillOffsetMemConfig_io_memData ),
       .io_outData( spillOffsetMem_io_outData ),
       .io_readEn( T728 ),
       .io_writeEn( spillOffsetMemConfig_io_memOutValid ),
       .io_readAddr( T727 ),
       .io_writeAddr( spillOffsetMemConfig_io_memAddr )
  );
  memConfig_1 loadSeqMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( loadSeqMemConfig_io_memAddr ),
       .io_memData( loadSeqMemConfig_io_memData ),
       .io_memOutValid( loadSeqMemConfig_io_memOutValid ),
       .io_rst( loadSeqMemConfig_io_rst )
  );
  memConfig_2 regLkupMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( regLkupMemConfig_io_memAddr ),
       .io_memData( regLkupMemConfig_io_memData ),
       .io_memOutValid( regLkupMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  memConfig_3 baseAddrMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( baseAddrMemConfig_io_memAddr ),
       .io_memData( baseAddrMemConfig_io_memData ),
       .io_memOutValid( baseAddrMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  memConfig_4 loopOffsetMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( loopOffsetMemConfig_io_memAddr ),
       .io_memData( loopOffsetMemConfig_io_memData ),
       .io_memOutValid( loopOffsetMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  memConfig_5 spillOffsetMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( spillOffsetMemConfig_io_memAddr ),
       .io_memData( spillOffsetMemConfig_io_memData ),
       .io_memOutValid( spillOffsetMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  fifo_2 lrRespFifo(.clk(clk), .reset(reset),
       .io_enqData( io_loadResp ),
       .io_deqData( lrRespFifo_io_deqData ),
       .io_enqRdy( lrRespFifo_io_enqRdy ),
       .io_deqRdy( lRespFifoDeq ),
       .io_enqValid( io_loadRespValid ),
       .io_deqValid( lrRespFifo_io_deqValid ),
       .io_rst( T716 )
  );
  fifo_3 lrReqFifo(.clk(clk), .reset(reset),
       .io_enqData( T768 ),
       .io_deqData( lrReqFifo_io_deqData ),
       .io_enqRdy( lrReqFifo_io_enqRdy ),
       .io_deqRdy( io_loadRqstRdy ),
       .io_enqValid( T238 ),
       .io_deqValid( lrReqFifo_io_deqValid ),
       .io_rst( T237 )
  );
  fifo_4 fifo(.clk(clk), .reset(reset),
       .io_enqData( T233 ),
       .io_deqData( fifo_io_deqData ),
       .io_enqRdy( fifo_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_0 ),
       .io_enqValid( T232 ),
       .io_deqValid( fifo_io_deqValid ),
       .io_rst( T231 )
  );
  fifo_4 fifo_1(.clk(clk), .reset(reset),
       .io_enqData( T227 ),
       .io_deqData( fifo_1_io_deqData ),
       .io_enqRdy( fifo_1_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_1 ),
       .io_enqValid( T226 ),
       .io_deqValid( fifo_1_io_deqValid ),
       .io_rst( T225 )
  );
  fifo_4 fifo_2(.clk(clk), .reset(reset),
       .io_enqData( T221 ),
       .io_deqData( fifo_2_io_deqData ),
       .io_enqRdy( fifo_2_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_2 ),
       .io_enqValid( T220 ),
       .io_deqValid( fifo_2_io_deqValid ),
       .io_rst( T219 )
  );
  fifo_4 fifo_3(.clk(clk), .reset(reset),
       .io_enqData( T215 ),
       .io_deqData( fifo_3_io_deqData ),
       .io_enqRdy( fifo_3_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_3 ),
       .io_enqValid( T214 ),
       .io_deqValid( fifo_3_io_deqValid ),
       .io_rst( T213 )
  );
  fifo_4 fifo_4(.clk(clk), .reset(reset),
       .io_enqData( T209 ),
       .io_deqData( fifo_4_io_deqData ),
       .io_enqRdy( fifo_4_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_4 ),
       .io_enqValid( T208 ),
       .io_deqValid( fifo_4_io_deqValid ),
       .io_rst( T207 )
  );
  fifo_4 fifo_5(.clk(clk), .reset(reset),
       .io_enqData( T203 ),
       .io_deqData( fifo_5_io_deqData ),
       .io_enqRdy( fifo_5_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_5 ),
       .io_enqValid( T202 ),
       .io_deqValid( fifo_5_io_deqValid ),
       .io_rst( T201 )
  );
  fifo_4 fifo_6(.clk(clk), .reset(reset),
       .io_enqData( T197 ),
       .io_deqData( fifo_6_io_deqData ),
       .io_enqRdy( fifo_6_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_6 ),
       .io_enqValid( T196 ),
       .io_deqValid( fifo_6_io_deqValid ),
       .io_rst( T195 )
  );
  fifo_4 fifo_7(.clk(clk), .reset(reset),
       .io_enqData( T188 ),
       .io_deqData( fifo_7_io_deqData ),
       .io_enqRdy( fifo_7_io_enqRdy ),
       .io_deqRdy( io_memBankRdy_7 ),
       .io_enqValid( T1 ),
       .io_deqValid( fifo_7_io_deqValid ),
       .io_rst( T0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      lRespDest <= 57'h0;
    end else if(T7) begin
      lRespDest <= regLookup;
    end
    if(reset) begin
      enqDoneReg <= 8'h0;
    end else if(T2) begin
      enqDoneReg <= T175;
    end else if(T174) begin
      enqDoneReg <= T166;
    end else if(T165) begin
      enqDoneReg <= T157;
    end else if(T156) begin
      enqDoneReg <= T148;
    end else if(T147) begin
      enqDoneReg <= T139;
    end else if(T138) begin
      enqDoneReg <= T130;
    end else if(T129) begin
      enqDoneReg <= T121;
    end else if(T120) begin
      enqDoneReg <= T112;
    end else begin
      enqDoneReg <= T18;
    end
    if(reset) begin
      lRespLkupValid <= 1'h0;
    end else if(T185) begin
      lRespLkupValid <= 1'h0;
    end else if(T7) begin
      lRespLkupValid <= 1'h1;
    end
    if(reset) begin
      lRespData <= 32'h0;
    end else if(T7) begin
      lRespData <= regLookupData;
    end
    if(reset) begin
      nextRqstValid <= 1'h0;
    end else if(T240) begin
      nextRqstValid <= 1'h0;
    end else if(seqInfoRegValid) begin
      nextRqstValid <= 1'h1;
    end
    if(reset) begin
      seqInfoRegValid <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      seqInfoRegValid <= 1'h0;
    end else if(seqInfoRegValid) begin
      seqInfoRegValid <= 1'h0;
    end else if(T247) begin
      seqInfoRegValid <= 1'h1;
    end
    nextRqst <= T769;
    if(reset) begin
      seqInfoReg <= 43'h0;
    end else if(T247) begin
      seqInfoReg <= loadSeqMem_io_outData;
    end
    if(reset) begin
      savedOffsets_0 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_0 <= 9'h0;
    end else if(T586) begin
      savedOffsets_0 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_1 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_1 <= 9'h0;
    end else if(T592) begin
      savedOffsets_1 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_2 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_2 <= 9'h0;
    end else if(T598) begin
      savedOffsets_2 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_3 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_3 <= 9'h0;
    end else if(T602) begin
      savedOffsets_3 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_4 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_4 <= 9'h0;
    end else if(T610) begin
      savedOffsets_4 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_5 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_5 <= 9'h0;
    end else if(T614) begin
      savedOffsets_5 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_6 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_6 <= 9'h0;
    end else if(T620) begin
      savedOffsets_6 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_7 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_7 <= 9'h0;
    end else if(T624) begin
      savedOffsets_7 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_8 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_8 <= 9'h0;
    end else if(T634) begin
      savedOffsets_8 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_9 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_9 <= 9'h0;
    end else if(T638) begin
      savedOffsets_9 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_10 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_10 <= 9'h0;
    end else if(T644) begin
      savedOffsets_10 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_11 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_11 <= 9'h0;
    end else if(T648) begin
      savedOffsets_11 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_12 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_12 <= 9'h0;
    end else if(T656) begin
      savedOffsets_12 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_13 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_13 <= 9'h0;
    end else if(T660) begin
      savedOffsets_13 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_14 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_14 <= 9'h0;
    end else if(T666) begin
      savedOffsets_14 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_15 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_15 <= 9'h0;
    end else if(T670) begin
      savedOffsets_15 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_16 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_16 <= 9'h0;
    end else if(T680) begin
      savedOffsets_16 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_17 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_17 <= 9'h0;
    end else if(T684) begin
      savedOffsets_17 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_18 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_18 <= 9'h0;
    end else if(T690) begin
      savedOffsets_18 <= savedOffsetsVal;
    end
    if(reset) begin
      savedOffsets_19 <= 9'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      savedOffsets_19 <= 9'h0;
    end else if(T694) begin
      savedOffsets_19 <= savedOffsetsVal;
    end
    if(reset) begin
      epilogueAfterSpill <= 1'h0;
    end else if(seqInfoRegValid) begin
      epilogueAfterSpill <= epilogueAfterSpillVal;
    end
    if(reset) begin
      spillEnd <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      spillEnd <= 1'h0;
    end else if(T247) begin
      spillEnd <= io_spillEnd;
    end
    if(reset) begin
      nextIterStart <= 1'h0;
    end else if(T247) begin
      nextIterStart <= io_nextIterStart;
    end
    if(reset) begin
      offsetUpdate_0 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_0 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_0 <= offsetUpdateVal_0;
    end
    if(reset) begin
      offsetUpdate_1 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_1 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_1 <= offsetUpdateVal_1;
    end
    if(reset) begin
      offsetUpdate_2 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_2 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_2 <= offsetUpdateVal_2;
    end
    if(reset) begin
      offsetUpdate_3 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_3 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_3 <= offsetUpdateVal_3;
    end
    if(reset) begin
      offsetUpdate_4 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_4 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_4 <= offsetUpdateVal_4;
    end
    if(reset) begin
      offsetUpdate_5 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_5 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_5 <= offsetUpdateVal_5;
    end
    if(reset) begin
      offsetUpdate_6 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_6 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_6 <= offsetUpdateVal_6;
    end
    if(reset) begin
      offsetUpdate_7 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_7 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_7 <= offsetUpdateVal_7;
    end
    if(reset) begin
      offsetUpdate_8 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_8 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_8 <= offsetUpdateVal_8;
    end
    if(reset) begin
      offsetUpdate_9 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_9 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_9 <= offsetUpdateVal_9;
    end
    if(reset) begin
      offsetUpdate_10 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_10 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_10 <= offsetUpdateVal_10;
    end
    if(reset) begin
      offsetUpdate_11 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_11 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_11 <= offsetUpdateVal_11;
    end
    if(reset) begin
      offsetUpdate_12 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_12 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_12 <= offsetUpdateVal_12;
    end
    if(reset) begin
      offsetUpdate_13 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_13 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_13 <= offsetUpdateVal_13;
    end
    if(reset) begin
      offsetUpdate_14 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_14 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_14 <= offsetUpdateVal_14;
    end
    if(reset) begin
      offsetUpdate_15 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_15 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_15 <= offsetUpdateVal_15;
    end
    if(reset) begin
      offsetUpdate_16 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_16 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_16 <= offsetUpdateVal_16;
    end
    if(reset) begin
      offsetUpdate_17 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_17 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_17 <= offsetUpdateVal_17;
    end
    if(reset) begin
      offsetUpdate_18 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_18 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_18 <= offsetUpdateVal_18;
    end
    if(reset) begin
      offsetUpdate_19 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      offsetUpdate_19 <= 1'h0;
    end else if(seqInfoRegValid) begin
      offsetUpdate_19 <= offsetUpdateVal_19;
    end
    if(reset) begin
      noCopyBaseAddr_0 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_0 <= 1'h0;
    end else if(T459) begin
      noCopyBaseAddr_0 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_1 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_1 <= 1'h0;
    end else if(T467) begin
      noCopyBaseAddr_1 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_2 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_2 <= 1'h0;
    end else if(T473) begin
      noCopyBaseAddr_2 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_3 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_3 <= 1'h0;
    end else if(T477) begin
      noCopyBaseAddr_3 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_4 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_4 <= 1'h0;
    end else if(T485) begin
      noCopyBaseAddr_4 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_5 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_5 <= 1'h0;
    end else if(T489) begin
      noCopyBaseAddr_5 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_6 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_6 <= 1'h0;
    end else if(T495) begin
      noCopyBaseAddr_6 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_7 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_7 <= 1'h0;
    end else if(T499) begin
      noCopyBaseAddr_7 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_8 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_8 <= 1'h0;
    end else if(T509) begin
      noCopyBaseAddr_8 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_9 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_9 <= 1'h0;
    end else if(T513) begin
      noCopyBaseAddr_9 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_10 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_10 <= 1'h0;
    end else if(T519) begin
      noCopyBaseAddr_10 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_11 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_11 <= 1'h0;
    end else if(T523) begin
      noCopyBaseAddr_11 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_12 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_12 <= 1'h0;
    end else if(T531) begin
      noCopyBaseAddr_12 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_13 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_13 <= 1'h0;
    end else if(T535) begin
      noCopyBaseAddr_13 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_14 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_14 <= 1'h0;
    end else if(T541) begin
      noCopyBaseAddr_14 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_15 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_15 <= 1'h0;
    end else if(T545) begin
      noCopyBaseAddr_15 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_16 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_16 <= 1'h0;
    end else if(T555) begin
      noCopyBaseAddr_16 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_17 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_17 <= 1'h0;
    end else if(T559) begin
      noCopyBaseAddr_17 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_18 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_18 <= 1'h0;
    end else if(T565) begin
      noCopyBaseAddr_18 <= 1'h1;
    end
    if(reset) begin
      noCopyBaseAddr_19 <= 1'h0;
    end else if(loadSeqMemConfig_io_rst) begin
      noCopyBaseAddr_19 <= 1'h0;
    end else if(T569) begin
      noCopyBaseAddr_19 <= 1'h1;
    end
    if(reset) begin
      lookupIndex <= 2'h0;
    end else if(T723) begin
      lookupIndex <= T738;
    end else if(T720) begin
      lookupIndex <= 2'h0;
    end
  end
endmodule

module loadSeq(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_loadRqst,
    output io_loadRqstValid,
    input  io_loadRqstRdy,
    input [37:0] io_loadResp,
    input  io_loadRespValid,
    output io_loadRespRdy,
    output[37:0] io_memBankEnq_7,
    output[37:0] io_memBankEnq_6,
    output[37:0] io_memBankEnq_5,
    output[37:0] io_memBankEnq_4,
    output[37:0] io_memBankEnq_3,
    output[37:0] io_memBankEnq_2,
    output[37:0] io_memBankEnq_1,
    output[37:0] io_memBankEnq_0,
    output io_memBankValid_7,
    output io_memBankValid_6,
    output io_memBankValid_5,
    output io_memBankValid_4,
    output io_memBankValid_3,
    output io_memBankValid_2,
    output io_memBankValid_1,
    output io_memBankValid_0,
    input  io_memBankRdy_7,
    input  io_memBankRdy_6,
    input  io_memBankRdy_5,
    input  io_memBankRdy_4,
    input  io_memBankRdy_3,
    input  io_memBankRdy_2,
    input  io_memBankRdy_1,
    input  io_memBankRdy_0
);

  wire loadCtrlClass_io_spillEnd;
  wire loadCtrlClass_io_nextIterStart;
  wire[8:0] loadCtrlClass_io_seqMemAddr;
  wire loadCtrlClass_io_seqMemAddrValid;
  wire[37:0] loadDPClass_io_memBankEnq_7;
  wire[37:0] loadDPClass_io_memBankEnq_6;
  wire[37:0] loadDPClass_io_memBankEnq_5;
  wire[37:0] loadDPClass_io_memBankEnq_4;
  wire[37:0] loadDPClass_io_memBankEnq_3;
  wire[37:0] loadDPClass_io_memBankEnq_2;
  wire[37:0] loadDPClass_io_memBankEnq_1;
  wire[37:0] loadDPClass_io_memBankEnq_0;
  wire loadDPClass_io_memBankValid_7;
  wire loadDPClass_io_memBankValid_6;
  wire loadDPClass_io_memBankValid_5;
  wire loadDPClass_io_memBankValid_4;
  wire loadDPClass_io_memBankValid_3;
  wire loadDPClass_io_memBankValid_2;
  wire loadDPClass_io_memBankValid_1;
  wire loadDPClass_io_memBankValid_0;
  wire[31:0] loadDPClass_io_loadRqst;
  wire loadDPClass_io_loadRqstValid;
  wire loadDPClass_io_loadRespRdy;
  wire loadDPClass_io_seqProceed;


  assign io_memBankValid_0 = loadDPClass_io_memBankValid_0;
  assign io_memBankValid_1 = loadDPClass_io_memBankValid_1;
  assign io_memBankValid_2 = loadDPClass_io_memBankValid_2;
  assign io_memBankValid_3 = loadDPClass_io_memBankValid_3;
  assign io_memBankValid_4 = loadDPClass_io_memBankValid_4;
  assign io_memBankValid_5 = loadDPClass_io_memBankValid_5;
  assign io_memBankValid_6 = loadDPClass_io_memBankValid_6;
  assign io_memBankValid_7 = loadDPClass_io_memBankValid_7;
  assign io_memBankEnq_0 = loadDPClass_io_memBankEnq_0;
  assign io_memBankEnq_1 = loadDPClass_io_memBankEnq_1;
  assign io_memBankEnq_2 = loadDPClass_io_memBankEnq_2;
  assign io_memBankEnq_3 = loadDPClass_io_memBankEnq_3;
  assign io_memBankEnq_4 = loadDPClass_io_memBankEnq_4;
  assign io_memBankEnq_5 = loadDPClass_io_memBankEnq_5;
  assign io_memBankEnq_6 = loadDPClass_io_memBankEnq_6;
  assign io_memBankEnq_7 = loadDPClass_io_memBankEnq_7;
  assign io_loadRespRdy = loadDPClass_io_loadRespRdy;
  assign io_loadRqstValid = loadDPClass_io_loadRqstValid;
  assign io_loadRqst = loadDPClass_io_loadRqst;
  loadSeqCtrl loadCtrlClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_spillEnd( loadCtrlClass_io_spillEnd ),
       .io_nextIterStart( loadCtrlClass_io_nextIterStart ),
       .io_seqMemAddr( loadCtrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( loadCtrlClass_io_seqMemAddrValid ),
       //.io_computeEnable(  )
       .io_seqProceed( loadDPClass_io_seqProceed )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign loadCtrlClass.io_seqMemAddrValid = {1{$random}};
// synthesis translate_on
`endif
  loadSeqDP loadDPClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_spillEnd( loadCtrlClass_io_spillEnd ),
       .io_nextIterStart( loadCtrlClass_io_nextIterStart ),
       .io_seqMemAddr( loadCtrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( loadCtrlClass_io_seqMemAddrValid ),
       .io_memBankEnq_7( loadDPClass_io_memBankEnq_7 ),
       .io_memBankEnq_6( loadDPClass_io_memBankEnq_6 ),
       .io_memBankEnq_5( loadDPClass_io_memBankEnq_5 ),
       .io_memBankEnq_4( loadDPClass_io_memBankEnq_4 ),
       .io_memBankEnq_3( loadDPClass_io_memBankEnq_3 ),
       .io_memBankEnq_2( loadDPClass_io_memBankEnq_2 ),
       .io_memBankEnq_1( loadDPClass_io_memBankEnq_1 ),
       .io_memBankEnq_0( loadDPClass_io_memBankEnq_0 ),
       .io_memBankValid_7( loadDPClass_io_memBankValid_7 ),
       .io_memBankValid_6( loadDPClass_io_memBankValid_6 ),
       .io_memBankValid_5( loadDPClass_io_memBankValid_5 ),
       .io_memBankValid_4( loadDPClass_io_memBankValid_4 ),
       .io_memBankValid_3( loadDPClass_io_memBankValid_3 ),
       .io_memBankValid_2( loadDPClass_io_memBankValid_2 ),
       .io_memBankValid_1( loadDPClass_io_memBankValid_1 ),
       .io_memBankValid_0( loadDPClass_io_memBankValid_0 ),
       .io_memBankRdy_7( io_memBankRdy_7 ),
       .io_memBankRdy_6( io_memBankRdy_6 ),
       .io_memBankRdy_5( io_memBankRdy_5 ),
       .io_memBankRdy_4( io_memBankRdy_4 ),
       .io_memBankRdy_3( io_memBankRdy_3 ),
       .io_memBankRdy_2( io_memBankRdy_2 ),
       .io_memBankRdy_1( io_memBankRdy_1 ),
       .io_memBankRdy_0( io_memBankRdy_0 ),
       .io_loadRqst( loadDPClass_io_loadRqst ),
       .io_loadRqstValid( loadDPClass_io_loadRqstValid ),
       .io_loadRqstRdy( io_loadRqstRdy ),
       .io_loadResp( io_loadResp ),
       .io_loadRespValid( io_loadRespValid ),
       .io_loadRespRdy( loadDPClass_io_loadRespRdy ),
       .io_seqProceed( loadDPClass_io_seqProceed )
  );
endmodule

module controllerConfigure_2(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_outConfig,
    output io_outValid,
    output io_computeCtrl,
    output io_computeCtrlValid
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  reg [31:0] inDataReg;
  wire[31:0] T30;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inDataReg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_computeCtrlValid = T0;
  assign T0 = T21 ? 1'h0 : T1;
  assign T1 = T18 ? 1'h1 : T2;
  assign T2 = T13 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : 1'h0;
  assign T4 = T11 & T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 2'h0;
  assign T7 = inDataReg[5'h1f:5'h1e];
  assign T30 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inDataReg;
  assign T9 = T10 == 1'h1;
  assign T10 = inDataReg[1'h0:1'h0];
  assign T11 = T12 == 1'h0;
  assign T12 = inDataReg[5'h1f:5'h1f];
  assign T13 = T11 & T14;
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h101;
  assign T16 = inDataReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T11 & T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T5 | T15;
  assign T21 = T11 ^ 1'h1;
  assign io_computeCtrl = T22;
  assign T22 = T21 ? 1'h0 : T23;
  assign T23 = T18 ? 1'h0 : T24;
  assign T24 = T13 ? 1'h0 : T25;
  assign T25 = T4 ? 1'h1 : 1'h0;
  assign io_outValid = T26;
  assign T26 = T21 ? 1'h0 : T27;
  assign T27 = T18 ? 1'h0 : T28;
  assign T28 = T13 ? 1'h1 : T29;
  assign T29 = T4 ? 1'h0 : 1'h0;
  assign io_outConfig = inDataReg;

  always @(posedge clk) begin
    if(reset) begin
      inDataReg <= 32'h0;
    end else if(io_inValid) begin
      inDataReg <= io_inConfig;
    end
  end
endmodule

module storeSeqCtrl(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output io_spillEnd,
    output io_nextIterStart,
    output[8:0] io_seqMemAddr,
    output io_seqMemAddrValid,
    input  io_seqProceed,
    output io_computeDone
);

  wire T0;
  reg  computeEnable;
  wire T130;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[514:0] lastAddr;
  wire[514:0] T131;
  wire[513:0] T7;
  wire[513:0] T132;
  reg [8:0] epilogueDepth;
  wire[8:0] T133;
  wire[8:0] T8;
  wire[8:0] T134;
  wire[6:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire[9:0] T22;
  wire[513:0] ssEnd;
  wire[513:0] T135;
  wire[8:0] T23;
  reg [8:0] steadyStateDepth;
  wire[8:0] T136;
  wire[9:0] T137;
  wire[9:0] T24;
  wire[9:0] T138;
  wire[9:0] T25;
  wire T26;
  reg [8:0] prologueDepth;
  wire[8:0] T139;
  wire[8:0] T27;
  wire[8:0] T140;
  wire[6:0] T28;
  wire startComputeValid;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire computeDone;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[514:0] T37;
  wire[514:0] T141;
  reg [511:0] seqMemAddr;
  wire[511:0] T142;
  wire[513:0] T143;
  wire[513:0] T38;
  wire[513:0] T39;
  wire[513:0] T144;
  wire[511:0] T40;
  wire[511:0] T41;
  wire[511:0] T42;
  wire T43;
  wire T44;
  wire nextRequest;
  wire T45;
  wire T46;
  wire T47;
  wire[511:0] T145;
  wire T48;
  wire T49;
  wire T50;
  reg [8:0] epilogueSpill;
  wire[8:0] T146;
  wire[9:0] T147;
  wire[9:0] T51;
  wire[9:0] T148;
  wire[9:0] T52;
  wire T53;
  wire[31:0] T54;
  reg [31:0] iterCount;
  wire[31:0] T149;
  wire[31:0] T55;
  wire[31:0] T150;
  wire[18:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire[2:0] T60;
  wire T61;
  reg [31:0] currentIter;
  wire[31:0] T151;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire T65;
  wire T66;
  wire[513:0] T67;
  wire[513:0] T152;
  wire T68;
  wire T69;
  wire[511:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[513:0] T77;
  wire[513:0] T153;
  wire T78;
  wire T79;
  wire[513:0] T154;
  wire[511:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[31:0] T91;
  wire T92;
  wire[514:0] T93;
  wire[514:0] T155;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[513:0] T101;
  wire[513:0] spillEndAddr;
  wire[513:0] T156;
  wire[8:0] T102;
  wire[513:0] T157;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire resetComputeValid;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[8:0] T158;
  wire[511:0] T117;
  wire[511:0] T118;
  wire T119;
  reg  nextIterStart;
  wire T159;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  reg  spillEnd;
  wire T160;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire storeCtrlConfigure_io_computeCtrl;
  wire storeCtrlConfigure_io_computeCtrlValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    computeEnable = {1{$random}};
    epilogueDepth = {1{$random}};
    steadyStateDepth = {1{$random}};
    prologueDepth = {1{$random}};
    seqMemAddr = {16{$random}};
    epilogueSpill = {1{$random}};
    iterCount = {1{$random}};
    currentIter = {1{$random}};
    nextIterStart = {1{$random}};
    spillEnd = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_computeDone = T0;
  assign T0 = computeEnable ^ 1'h1;
  assign T130 = reset ? 1'h0 : T1;
  assign T1 = T113 ? 1'h0 : T2;
  assign T2 = T110 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : computeEnable;
  assign T4 = T32 & T5;
  assign T5 = startComputeValid & T6;
  assign T6 = lastAddr != 515'h0;
  assign lastAddr = T131;
  assign T131 = {1'h0, T7};
  assign T7 = ssEnd + T132;
  assign T132 = {505'h0, epilogueDepth};
  assign T133 = reset ? 9'h0 : T8;
  assign T8 = T10 ? T134 : epilogueDepth;
  assign T134 = {2'h0, T9};
  assign T9 = io_inConfig[3'h6:1'h0];
  assign T10 = T17 & T11;
  assign T11 = T14 & T12;
  assign T12 = T13 == 1'h1;
  assign T13 = io_inConfig[5'h11:5'h11];
  assign T14 = T15 ^ 1'h1;
  assign T15 = T16 == 1'h0;
  assign T16 = io_inConfig[5'h11:5'h11];
  assign T17 = T20 & T18;
  assign T18 = T19 == 3'h0;
  assign T19 = io_inConfig[5'h15:5'h13];
  assign T20 = io_inValid & T21;
  assign T21 = T22 == 10'h103;
  assign T22 = io_inConfig[5'h1f:5'h16];
  assign ssEnd = T135;
  assign T135 = {505'h0, T23};
  assign T23 = prologueDepth + steadyStateDepth;
  assign T136 = T137[4'h8:1'h0];
  assign T137 = reset ? 10'h0 : T24;
  assign T24 = T26 ? T25 : T138;
  assign T138 = {1'h0, steadyStateDepth};
  assign T25 = io_inConfig[5'h10:3'h7];
  assign T26 = T17 & T15;
  assign T139 = reset ? 9'h0 : T27;
  assign T27 = T26 ? T140 : prologueDepth;
  assign T140 = {2'h0, T28};
  assign T28 = io_inConfig[3'h6:1'h0];
  assign startComputeValid = T29;
  assign T29 = T31 ? 1'h0 : T30;
  assign T30 = storeCtrlConfigure_io_computeCtrlValid & storeCtrlConfigure_io_computeCtrl;
  assign T31 = storeCtrlConfigure_io_computeCtrlValid ^ 1'h1;
  assign T32 = T106 | computeDone;
  assign computeDone = T33;
  assign T33 = T103 ? T98 : T34;
  assign T34 = T94 ? T89 : T35;
  assign T35 = T84 ? T36 : 1'h0;
  assign T36 = T141 == T37;
  assign T37 = lastAddr - 515'h1;
  assign T141 = {3'h0, seqMemAddr};
  assign T142 = T143[9'h1ff:1'h0];
  assign T143 = reset ? 514'h0 : T38;
  assign T38 = T81 ? T154 : T39;
  assign T39 = T73 ? ssEnd : T144;
  assign T144 = {2'h0, T40};
  assign T40 = T71 ? T70 : T41;
  assign T41 = T48 ? T145 : T42;
  assign T42 = T43 ? 512'h0 : seqMemAddr;
  assign T43 = T44 & startComputeValid;
  assign T44 = startComputeValid | nextRequest;
  assign nextRequest = T45;
  assign T45 = T47 ? 1'h0 : T46;
  assign T46 = io_seqProceed & computeEnable;
  assign T47 = T46 ^ 1'h1;
  assign T145 = {503'h0, prologueDepth};
  assign T48 = T65 & T49;
  assign T49 = T53 | T50;
  assign T50 = epilogueSpill != 9'h0;
  assign T146 = T147[4'h8:1'h0];
  assign T147 = reset ? 10'h0 : T51;
  assign T51 = T10 ? T52 : T148;
  assign T148 = {1'h0, epilogueSpill};
  assign T52 = io_inConfig[5'h10:3'h7];
  assign T53 = currentIter < T54;
  assign T54 = iterCount - 32'h1;
  assign T149 = reset ? 32'h0 : T55;
  assign T55 = T57 ? T150 : iterCount;
  assign T150 = {13'h0, T56};
  assign T56 = io_inConfig[5'h12:1'h0];
  assign T57 = T20 & T58;
  assign T58 = T61 & T59;
  assign T59 = T60 == 3'h1;
  assign T60 = io_inConfig[5'h15:5'h13];
  assign T61 = T18 ^ 1'h1;
  assign T151 = reset ? 32'h0 : T62;
  assign T62 = T48 ? T64 : T63;
  assign T63 = T43 ? 32'h0 : currentIter;
  assign T64 = currentIter + 32'h1;
  assign T65 = T68 & T66;
  assign T66 = T152 == T67;
  assign T67 = ssEnd - 514'h1;
  assign T152 = {2'h0, seqMemAddr};
  assign T68 = T44 & T69;
  assign T69 = startComputeValid ^ 1'h1;
  assign T70 = seqMemAddr + 512'h1;
  assign T71 = T65 & T72;
  assign T72 = T49 ^ 1'h1;
  assign T73 = T68 & T74;
  assign T74 = T79 & T75;
  assign T75 = T78 & T76;
  assign T76 = T153 == T77;
  assign T77 = ssEnd - 514'h1;
  assign T153 = {2'h0, seqMemAddr};
  assign T78 = currentIter == iterCount;
  assign T79 = T66 ^ 1'h1;
  assign T154 = {2'h0, T80};
  assign T80 = seqMemAddr + 512'h1;
  assign T81 = T68 & T82;
  assign T82 = T83 ^ 1'h1;
  assign T83 = T66 | T75;
  assign T84 = T88 & T85;
  assign T85 = T87 & T86;
  assign T86 = steadyStateDepth == 9'h1;
  assign T87 = epilogueDepth != 9'h0;
  assign T88 = computeEnable & nextRequest;
  assign T89 = T92 & T90;
  assign T90 = T91 == iterCount;
  assign T91 = currentIter + 32'h1;
  assign T92 = T155 == T93;
  assign T93 = lastAddr - 515'h1;
  assign T155 = {3'h0, seqMemAddr};
  assign T94 = T88 & T95;
  assign T95 = T97 & T96;
  assign T96 = epilogueSpill == 9'h0;
  assign T97 = T85 ^ 1'h1;
  assign T98 = T100 & T99;
  assign T99 = currentIter == iterCount;
  assign T100 = T157 == T101;
  assign T101 = spillEndAddr - 514'h1;
  assign spillEndAddr = T156;
  assign T156 = {505'h0, T102};
  assign T102 = prologueDepth + epilogueSpill;
  assign T157 = {2'h0, seqMemAddr};
  assign T103 = T88 & T104;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T85 | T96;
  assign T106 = startComputeValid | resetComputeValid;
  assign resetComputeValid = T107;
  assign T107 = T31 ? 1'h0 : T108;
  assign T108 = storeCtrlConfigure_io_computeCtrlValid & T109;
  assign T109 = storeCtrlConfigure_io_computeCtrl ^ 1'h1;
  assign T110 = T32 & T111;
  assign T111 = T112 & resetComputeValid;
  assign T112 = T5 ^ 1'h1;
  assign T113 = T32 & T114;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T5 | resetComputeValid;
  assign io_seqMemAddrValid = T116;
  assign T116 = T46 ? 1'h1 : 1'h0;
  assign io_seqMemAddr = T158;
  assign T158 = T117[4'h8:1'h0];
  assign T117 = T46 ? seqMemAddr : T118;
  assign T118 = T44 ? seqMemAddr : seqMemAddr;
  assign io_nextIterStart = T119;
  assign T119 = T46 ? nextIterStart : nextIterStart;
  assign T159 = reset ? 1'h0 : T120;
  assign T120 = T81 ? 1'h0 : T121;
  assign T121 = T73 ? 1'h0 : T122;
  assign T122 = T71 ? 1'h0 : T123;
  assign T123 = T48 ? 1'h1 : T124;
  assign T124 = T43 ? 1'h0 : nextIterStart;
  assign io_spillEnd = T125;
  assign T125 = T46 ? spillEnd : spillEnd;
  assign T160 = reset ? 1'h0 : T126;
  assign T126 = T81 ? 1'h0 : T127;
  assign T127 = T73 ? 1'h1 : T128;
  assign T128 = T65 ? 1'h0 : T129;
  assign T129 = T43 ? 1'h0 : spillEnd;
  controllerConfigure_2 storeCtrlConfigure(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       //.io_outConfig(  )
       //.io_outValid(  )
       .io_computeCtrl( storeCtrlConfigure_io_computeCtrl ),
       .io_computeCtrlValid( storeCtrlConfigure_io_computeCtrlValid )
  );

  always @(posedge clk) begin
    if(reset) begin
      computeEnable <= 1'h0;
    end else if(T113) begin
      computeEnable <= 1'h0;
    end else if(T110) begin
      computeEnable <= 1'h0;
    end else if(T4) begin
      computeEnable <= 1'h1;
    end
    if(reset) begin
      epilogueDepth <= 9'h0;
    end else if(T10) begin
      epilogueDepth <= T134;
    end
    steadyStateDepth <= T136;
    if(reset) begin
      prologueDepth <= 9'h0;
    end else if(T26) begin
      prologueDepth <= T140;
    end
    seqMemAddr <= T142;
    epilogueSpill <= T146;
    if(reset) begin
      iterCount <= 32'h0;
    end else if(T57) begin
      iterCount <= T150;
    end
    if(reset) begin
      currentIter <= 32'h0;
    end else if(T48) begin
      currentIter <= T64;
    end else if(T43) begin
      currentIter <= 32'h0;
    end
    if(reset) begin
      nextIterStart <= 1'h0;
    end else if(T81) begin
      nextIterStart <= 1'h0;
    end else if(T73) begin
      nextIterStart <= 1'h0;
    end else if(T71) begin
      nextIterStart <= 1'h0;
    end else if(T48) begin
      nextIterStart <= 1'h1;
    end else if(T43) begin
      nextIterStart <= 1'h0;
    end
    if(reset) begin
      spillEnd <= 1'h0;
    end else if(T81) begin
      spillEnd <= 1'h0;
    end else if(T73) begin
      spillEnd <= 1'h1;
    end else if(T65) begin
      spillEnd <= 1'h0;
    end else if(T43) begin
      spillEnd <= 1'h0;
    end
  end
endmodule

module memConfig_6(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[8:0] io_memAddr,
    output[42:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[5:0] T94;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[5:0] T95;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[5:0] T96;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[5:0] T97;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[42:0] T98;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T99;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T100;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[8:0] T87;
  reg [8:0] memAddr;
  wire[8:0] T101;
  wire[8:0] T88;
  wire[8:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T94 == 6'h20;
  assign T94 = {1'h0, T58};
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T95 == 6'h20;
  assign T95 = {1'h0, T63};
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T96 == 6'h20;
  assign T96 = {1'h0, T68};
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T97 == 6'h20;
  assign T97 = {1'h0, T73};
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T98;
  assign T98 = T76[6'h2a:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T99 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T100 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 9'h0;
  assign T101 = reset ? 9'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 9'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 9'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_7(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[5:0] T94;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[5:0] T95;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[5:0] T96;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[5:0] T97;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T98;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T99;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T100;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T101;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T94 == 6'h21;
  assign T94 = {1'h0, T58};
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T95 == 6'h21;
  assign T95 = {1'h0, T63};
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T96 == 6'h21;
  assign T96 = {1'h0, T68};
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T97 == 6'h21;
  assign T97 = {1'h0, T73};
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T98;
  assign T98 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T99 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T100 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T101 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_8(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[5:0] T94;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[5:0] T95;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[5:0] T96;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[5:0] T97;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T98;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T99;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T100;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T101;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T94 == 6'h22;
  assign T94 = {1'h0, T58};
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T95 == 6'h22;
  assign T95 = {1'h0, T63};
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T96 == 6'h22;
  assign T96 = {1'h0, T68};
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T97 == 6'h22;
  assign T97 = {1'h0, T73};
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T98;
  assign T98 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T99 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T100 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T101 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module memConfig_9(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[4:0] io_memAddr,
    output[31:0] io_memData,
    output io_memOutValid,
    output io_rst
);

  wire T0;
  wire startCompute;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [31:0] inConfigReg;
  wire[31:0] T90;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[9:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[9:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  memOutValid;
  wire T91;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg  iterCnt;
  wire T92;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  memTypeMatch;
  wire T93;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[5:0] T94;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[5:0] T95;
  wire[4:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[5:0] T96;
  wire[4:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[5:0] T97;
  wire[4:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T98;
  wire[61:0] T76;
  wire[61:0] T77;
  reg [30:0] memData_0;
  wire[30:0] T99;
  wire[30:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  reg [30:0] memData_1;
  wire[30:0] T100;
  wire[30:0] T84;
  wire T85;
  wire T86;
  wire[4:0] T87;
  reg [4:0] memAddr;
  wire[4:0] T101;
  wire[4:0] T88;
  wire[4:0] T89;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    inConfigReg = {1{$random}};
    memOutValid = {1{$random}};
    iterCnt = {1{$random}};
    memTypeMatch = {1{$random}};
    memData_0 = {1{$random}};
    memData_1 = {1{$random}};
    memAddr = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_rst = T0;
  assign T0 = startCompute ? 1'h1 : 1'h0;
  assign startCompute = T1;
  assign T1 = T28 ? 1'h0 : T2;
  assign T2 = T23 ? 1'h0 : T3;
  assign T3 = T18 ? 1'h0 : T4;
  assign T4 = T14 ? 1'h0 : T5;
  assign T5 = T9 & T6;
  assign T6 = T7 == 1'h1;
  assign T7 = inConfigReg[1'h0:1'h0];
  assign T90 = reset ? 32'h0 : T8;
  assign T8 = io_inValid ? io_inConfig : inConfigReg;
  assign T9 = T12 & T10;
  assign T10 = T11 == 2'h0;
  assign T11 = inConfigReg[5'h1e:5'h1d];
  assign T12 = T13 == 1'h0;
  assign T13 = inConfigReg[5'h1f:5'h1f];
  assign T14 = T17 & T15;
  assign T15 = T16 == 10'h100;
  assign T16 = inConfigReg[5'h1f:5'h16];
  assign T17 = T5 ^ 1'h1;
  assign T18 = T21 & T19;
  assign T19 = T20 == 10'h103;
  assign T20 = inConfigReg[5'h1f:5'h16];
  assign T21 = T22 ^ 1'h1;
  assign T22 = T5 | T15;
  assign T23 = T26 & T24;
  assign T24 = T25 == 10'h101;
  assign T25 = inConfigReg[5'h1f:5'h16];
  assign T26 = T27 ^ 1'h1;
  assign T27 = T22 | T19;
  assign T28 = T31 & T29;
  assign T29 = T30 == 10'h100;
  assign T30 = inConfigReg[5'h1f:5'h16];
  assign T31 = T32 ^ 1'h1;
  assign T32 = T27 | T24;
  assign io_memOutValid = T33;
  assign T33 = memOutValid ? 1'h1 : 1'h0;
  assign T91 = reset ? 1'h0 : T34;
  assign T34 = memOutValid ? 1'h0 : T35;
  assign T35 = T36 ? 1'h1 : memOutValid;
  assign T36 = T45 & T37;
  assign T37 = T44 & T38;
  assign T38 = iterCnt == 1'h1;
  assign T92 = reset ? 1'h0 : T39;
  assign T39 = T36 ? 1'h0 : T40;
  assign T40 = T42 ? T41 : iterCnt;
  assign T41 = iterCnt + 1'h1;
  assign T42 = T45 & T43;
  assign T43 = iterCnt < 1'h1;
  assign T44 = T43 ^ 1'h1;
  assign T45 = memTypeMatch & T46;
  assign T46 = T47 == 1'h1;
  assign T47 = inConfigReg[5'h1f:5'h1f];
  assign T93 = reset ? 1'h0 : T48;
  assign T48 = T74 ? 1'h0 : T49;
  assign T49 = T71 ? 1'h1 : T50;
  assign T50 = T69 ? 1'h0 : T51;
  assign T51 = T66 ? 1'h1 : T52;
  assign T52 = T64 ? 1'h0 : T53;
  assign T53 = T61 ? 1'h1 : T54;
  assign T54 = T59 ? 1'h0 : T55;
  assign T55 = T56 ? 1'h1 : memTypeMatch;
  assign T56 = T14 & T57;
  assign T57 = T94 == 6'h23;
  assign T94 = {1'h0, T58};
  assign T58 = inConfigReg[5'h17:5'h13];
  assign T59 = T14 & T60;
  assign T60 = T57 ^ 1'h1;
  assign T61 = T18 & T62;
  assign T62 = T95 == 6'h23;
  assign T95 = {1'h0, T63};
  assign T63 = inConfigReg[5'h17:5'h13];
  assign T64 = T18 & T65;
  assign T65 = T62 ^ 1'h1;
  assign T66 = T23 & T67;
  assign T67 = T96 == 6'h23;
  assign T96 = {1'h0, T68};
  assign T68 = inConfigReg[5'h17:5'h13];
  assign T69 = T23 & T70;
  assign T70 = T67 ^ 1'h1;
  assign T71 = T28 & T72;
  assign T72 = T97 == 6'h23;
  assign T97 = {1'h0, T73};
  assign T73 = inConfigReg[5'h17:5'h13];
  assign T74 = T28 & T75;
  assign T75 = T72 ^ 1'h1;
  assign io_memData = T98;
  assign T98 = T76[5'h1f:1'h0];
  assign T76 = memOutValid ? T77 : 62'h0;
  assign T77 = {memData_1, memData_0};
  assign T99 = reset ? 31'h0 : T78;
  assign T78 = T80 ? T79 : memData_0;
  assign T79 = inConfigReg[5'h1e:1'h0];
  assign T80 = T45 & T81;
  assign T81 = T82[1'h0:1'h0];
  assign T82 = 1'h1 << T83;
  assign T83 = iterCnt;
  assign T100 = reset ? 31'h0 : T84;
  assign T84 = T85 ? T79 : memData_1;
  assign T85 = T45 & T86;
  assign T86 = T82[1'h1:1'h1];
  assign io_memAddr = T87;
  assign T87 = memOutValid ? memAddr : 5'h0;
  assign T101 = reset ? 5'h0 : T88;
  assign T88 = memOutValid ? T89 : memAddr;
  assign T89 = memAddr + 5'h1;

  always @(posedge clk) begin
    if(reset) begin
      inConfigReg <= 32'h0;
    end else if(io_inValid) begin
      inConfigReg <= io_inConfig;
    end
    if(reset) begin
      memOutValid <= 1'h0;
    end else if(memOutValid) begin
      memOutValid <= 1'h0;
    end else if(T36) begin
      memOutValid <= 1'h1;
    end
    if(reset) begin
      iterCnt <= 1'h0;
    end else if(T36) begin
      iterCnt <= 1'h0;
    end else if(T42) begin
      iterCnt <= T41;
    end
    if(reset) begin
      memTypeMatch <= 1'h0;
    end else if(T74) begin
      memTypeMatch <= 1'h0;
    end else if(T71) begin
      memTypeMatch <= 1'h1;
    end else if(T69) begin
      memTypeMatch <= 1'h0;
    end else if(T66) begin
      memTypeMatch <= 1'h1;
    end else if(T64) begin
      memTypeMatch <= 1'h0;
    end else if(T61) begin
      memTypeMatch <= 1'h1;
    end else if(T59) begin
      memTypeMatch <= 1'h0;
    end else if(T56) begin
      memTypeMatch <= 1'h1;
    end
    if(reset) begin
      memData_0 <= 31'h0;
    end else if(T80) begin
      memData_0 <= T79;
    end
    if(reset) begin
      memData_1 <= 31'h0;
    end else if(T85) begin
      memData_1 <= T79;
    end
    if(reset) begin
      memAddr <= 5'h0;
    end else if(memOutValid) begin
      memAddr <= T89;
    end
  end
endmodule

module fifo_5(input clk, input reset,
    input [63:0] io_enqData,
    output[63:0] io_deqData,
    output io_enqRdy,
    input  io_deqRdy,
    input  io_enqValid,
    output io_deqValid,
    input  io_rst
);

  wire T0;
  wire isEmpty;
  wire T1;
  reg [2:0] deqPtr;
  wire[2:0] T21;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] deqPtrInc;
  wire[2:0] T4;
  wire doDeq;
  wire T5;
  reg [2:0] enqPtr;
  wire[2:0] T22;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] enqPtrInc;
  wire[2:0] T8;
  wire doEnq;
  wire T9;
  wire T10;
  reg  isFull;
  wire T23;
  wire T11;
  wire isFullNext;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[63:0] T19;
  reg [63:0] fifoMem [7:0];
  wire[63:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deqPtr = {1{$random}};
    enqPtr = {1{$random}};
    isFull = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      fifoMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_deqValid = T0;
  assign T0 = isEmpty ^ 1'h1;
  assign isEmpty = T10 & T1;
  assign T1 = enqPtr == deqPtr;
  assign T21 = reset ? 3'h0 : T2;
  assign T2 = io_rst ? 3'h0 : T3;
  assign T3 = doDeq ? deqPtrInc : deqPtr;
  assign deqPtrInc = T4 % 4'h8;
  assign T4 = deqPtr + 3'h1;
  assign doDeq = T5;
  assign T5 = io_deqValid & io_deqRdy;
  assign T22 = reset ? 3'h0 : T6;
  assign T6 = io_rst ? 3'h0 : T7;
  assign T7 = doEnq ? enqPtrInc : enqPtr;
  assign enqPtrInc = T8 % 4'h8;
  assign T8 = enqPtr + 3'h1;
  assign doEnq = T9;
  assign T9 = io_enqRdy & io_enqValid;
  assign T10 = isFull ^ 1'h1;
  assign T23 = reset ? 1'h0 : T11;
  assign T11 = io_rst ? 1'h0 : isFullNext;
  assign isFullNext = T14 ? 1'h1 : T12;
  assign T12 = T13 ? 1'h0 : isFull;
  assign T13 = doDeq & isFull;
  assign T14 = T16 & T15;
  assign T15 = enqPtrInc == deqPtr;
  assign T16 = doEnq & T17;
  assign T17 = ~ doDeq;
  assign io_enqRdy = T18;
  assign T18 = isFull ^ 1'h1;
  assign io_deqData = T19;
  assign T19 = fifoMem[deqPtr];

  always @(posedge clk) begin
    if(reset) begin
      deqPtr <= 3'h0;
    end else if(io_rst) begin
      deqPtr <= 3'h0;
    end else if(doDeq) begin
      deqPtr <= deqPtrInc;
    end
    if(reset) begin
      enqPtr <= 3'h0;
    end else if(io_rst) begin
      enqPtr <= 3'h0;
    end else if(doEnq) begin
      enqPtr <= enqPtrInc;
    end
    if(reset) begin
      isFull <= 1'h0;
    end else if(io_rst) begin
      isFull <= 1'h0;
    end else if(T14) begin
      isFull <= 1'h1;
    end else if(T13) begin
      isFull <= 1'h0;
    end
    if (doEnq)
      fifoMem[enqPtr] <= io_enqData;
  end
endmodule

module storeSeqDP(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input  io_spillEnd,
    input  io_nextIterStart,
    input [8:0] io_seqMemAddr,
    input  io_seqMemAddrValid,
    output[63:0] io_storeMemData,
    output io_storeMemValid,
    input  io_storeMemRdy,
    output io_seqProceed,
    input [31:0] io_fabOutToStore_19,
    input [31:0] io_fabOutToStore_18,
    input [31:0] io_fabOutToStore_17,
    input [31:0] io_fabOutToStore_16,
    input [31:0] io_fabOutToStore_15,
    input [31:0] io_fabOutToStore_14,
    input [31:0] io_fabOutToStore_13,
    input [31:0] io_fabOutToStore_12,
    input [31:0] io_fabOutToStore_11,
    input [31:0] io_fabOutToStore_10,
    input [31:0] io_fabOutToStore_9,
    input [31:0] io_fabOutToStore_8,
    input [31:0] io_fabOutToStore_7,
    input [31:0] io_fabOutToStore_6,
    input [31:0] io_fabOutToStore_5,
    input [31:0] io_fabOutToStore_4,
    input [31:0] io_fabOutToStore_3,
    input [31:0] io_fabOutToStore_2,
    input [31:0] io_fabOutToStore_1,
    input [31:0] io_fabOutToStore_0,
    input  io_fabOutToStoreValid_19,
    input  io_fabOutToStoreValid_18,
    input  io_fabOutToStoreValid_17,
    input  io_fabOutToStoreValid_16,
    input  io_fabOutToStoreValid_15,
    input  io_fabOutToStoreValid_14,
    input  io_fabOutToStoreValid_13,
    input  io_fabOutToStoreValid_12,
    input  io_fabOutToStoreValid_11,
    input  io_fabOutToStoreValid_10,
    input  io_fabOutToStoreValid_9,
    input  io_fabOutToStoreValid_8,
    input  io_fabOutToStoreValid_7,
    input  io_fabOutToStoreValid_6,
    input  io_fabOutToStoreValid_5,
    input  io_fabOutToStoreValid_4,
    input  io_fabOutToStoreValid_3,
    input  io_fabOutToStoreValid_2,
    input  io_fabOutToStoreValid_1,
    input  io_fabOutToStoreValid_0,
    output io_computeDone,
    input  io_computeDoneCtrl
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg  portSel_0;
  wire T881;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[31:0] T46;
  wire[4:0] T47;
  wire[4:0] portID;
  wire[4:0] T48;
  wire[4:0] T49;
  reg [42:0] nextSeq;
  wire[42:0] T882;
  wire[42:0] T50;
  wire T51;
  reg  nextSeqValid;
  wire T883;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  reg  firstReqDone;
  wire T884;
  wire T57;
  wire T58;
  wire getNextReq;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg  portSel_1;
  wire T885;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  portSel_2;
  wire T886;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  reg  portSel_3;
  wire T887;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  reg  portSel_4;
  wire T888;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  reg  portSel_5;
  wire T889;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  reg  portSel_6;
  wire T890;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  reg  portSel_7;
  wire T891;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  reg  portSel_8;
  wire T892;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  reg  portSel_9;
  wire T893;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  reg  portSel_10;
  wire T894;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  reg  portSel_11;
  wire T895;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  reg  portSel_12;
  wire T896;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  reg  portSel_13;
  wire T897;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  portSel_14;
  wire T898;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg  portSel_15;
  wire T899;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  reg  portSel_16;
  wire T900;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  reg  portSel_17;
  wire T901;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  reg  portSel_18;
  wire T902;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  reg  portSel_19;
  wire T903;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire[63:0] T233;
  wire[63:0] T234;
  wire[63:0] T235;
  wire[63:0] T236;
  wire[63:0] T237;
  wire[63:0] T238;
  wire[63:0] T239;
  wire[63:0] T240;
  wire[63:0] T241;
  wire[63:0] T242;
  wire[63:0] T243;
  wire[63:0] T244;
  wire[63:0] T245;
  wire[63:0] T246;
  wire[63:0] T247;
  wire[63:0] T248;
  wire[63:0] T249;
  wire[63:0] T250;
  wire[63:0] T251;
  wire[63:0] T252;
  wire[63:0] T253;
  wire[63:0] T254;
  wire[63:0] T255;
  wire[63:0] T256;
  wire[63:0] T257;
  wire[63:0] T258;
  wire[63:0] T259;
  wire[63:0] T260;
  wire[63:0] T261;
  wire[63:0] T262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire[63:0] T265;
  wire[63:0] T266;
  wire[63:0] T267;
  wire[63:0] T268;
  wire[63:0] T269;
  wire[63:0] T270;
  wire[63:0] T271;
  wire[63:0] T272;
  wire[31:0] storeReqData;
  wire[31:0] T273;
  wire[31:0] T274;
  wire[31:0] T275;
  wire[31:0] T276;
  wire[31:0] T277;
  wire[31:0] T278;
  wire[31:0] T279;
  wire[31:0] T280;
  wire[31:0] T281;
  wire[31:0] T282;
  wire[31:0] T283;
  wire[31:0] T284;
  wire[31:0] T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire[31:0] T288;
  wire[31:0] T289;
  wire[31:0] T290;
  wire[31:0] T291;
  wire[31:0] T292;
  wire[31:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[31:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[31:0] T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] storeReqAddr;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  wire[31:0] T322;
  wire[31:0] T323;
  wire[31:0] T324;
  wire[31:0] T325;
  wire[31:0] T326;
  wire[31:0] T327;
  wire[31:0] T328;
  wire[31:0] T329;
  wire[31:0] T330;
  wire[31:0] T331;
  wire[31:0] T332;
  wire[31:0] T333;
  wire[31:0] T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  wire[31:0] T344;
  wire[31:0] T345;
  wire[31:0] T346;
  wire[31:0] T347;
  wire[31:0] T348;
  wire[31:0] T349;
  wire[31:0] T350;
  wire[31:0] T351;
  wire[31:0] T352;
  reg [31:0] storeMemAddr;
  wire[31:0] T904;
  wire[31:0] T353;
  wire[31:0] T354;
  wire[31:0] offsetAddr;
  wire[31:0] T355;
  wire[31:0] T356;
  wire[31:0] T905;
  wire T357;
  wire T358;
  wire T359;
  wire[4:0] T360;
  wire[4:0] T361;
  wire[4:0] addrLkupIndex;
  wire[4:0] T362;
  wire[4:0] T363;
  wire T364;
  wire[8:0] savedOffsetsVal;
  wire[8:0] T906;
  wire[31:0] T365;
  wire[31:0] T366;
  wire[31:0] T367;
  wire[31:0] T368;
  wire[31:0] T369;
  wire[31:0] T370;
  wire[31:0] T371;
  wire[31:0] spillLkup;
  wire[31:0] T372;
  wire[31:0] T907;
  wire[8:0] T672;
  wire[8:0] T673;
  wire[8:0] T674;
  wire[8:0] T675;
  wire[8:0] T676;
  reg [8:0] savedOffsets_0;
  wire[8:0] T908;
  wire[8:0] T677;
  wire[8:0] T678;
  wire T679;
  wire T680;
  wire[31:0] T681;
  wire[4:0] T682;
  reg [8:0] savedOffsets_1;
  wire[8:0] T909;
  wire[8:0] T683;
  wire[8:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[8:0] T688;
  reg [8:0] savedOffsets_2;
  wire[8:0] T910;
  wire[8:0] T689;
  wire[8:0] T690;
  wire T691;
  wire T692;
  reg [8:0] savedOffsets_3;
  wire[8:0] T911;
  wire[8:0] T693;
  wire[8:0] T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire[8:0] T699;
  wire[8:0] T700;
  reg [8:0] savedOffsets_4;
  wire[8:0] T912;
  wire[8:0] T701;
  wire[8:0] T702;
  wire T703;
  wire T704;
  reg [8:0] savedOffsets_5;
  wire[8:0] T913;
  wire[8:0] T705;
  wire[8:0] T706;
  wire T707;
  wire T708;
  wire T709;
  wire[8:0] T710;
  reg [8:0] savedOffsets_6;
  wire[8:0] T914;
  wire[8:0] T711;
  wire[8:0] T712;
  wire T713;
  wire T714;
  reg [8:0] savedOffsets_7;
  wire[8:0] T915;
  wire[8:0] T715;
  wire[8:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire[8:0] T722;
  wire[8:0] T723;
  wire[8:0] T724;
  reg [8:0] savedOffsets_8;
  wire[8:0] T916;
  wire[8:0] T725;
  wire[8:0] T726;
  wire T727;
  wire T728;
  reg [8:0] savedOffsets_9;
  wire[8:0] T917;
  wire[8:0] T729;
  wire[8:0] T730;
  wire T731;
  wire T732;
  wire T733;
  wire[8:0] T734;
  reg [8:0] savedOffsets_10;
  wire[8:0] T918;
  wire[8:0] T735;
  wire[8:0] T736;
  wire T737;
  wire T738;
  reg [8:0] savedOffsets_11;
  wire[8:0] T919;
  wire[8:0] T739;
  wire[8:0] T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire[8:0] T745;
  wire[8:0] T746;
  reg [8:0] savedOffsets_12;
  wire[8:0] T920;
  wire[8:0] T747;
  wire[8:0] T748;
  wire T749;
  wire T750;
  reg [8:0] savedOffsets_13;
  wire[8:0] T921;
  wire[8:0] T751;
  wire[8:0] T752;
  wire T753;
  wire T754;
  wire T755;
  wire[8:0] T756;
  reg [8:0] savedOffsets_14;
  wire[8:0] T922;
  wire[8:0] T757;
  wire[8:0] T758;
  wire T759;
  wire T760;
  reg [8:0] savedOffsets_15;
  wire[8:0] T923;
  wire[8:0] T761;
  wire[8:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire T768;
  wire[8:0] T769;
  wire[8:0] T770;
  reg [8:0] savedOffsets_16;
  wire[8:0] T924;
  wire[8:0] T771;
  wire[8:0] T772;
  wire T773;
  wire T774;
  reg [8:0] savedOffsets_17;
  wire[8:0] T925;
  wire[8:0] T775;
  wire[8:0] T776;
  wire T777;
  wire T778;
  wire T779;
  wire[8:0] T780;
  reg [8:0] savedOffsets_18;
  wire[8:0] T926;
  wire[8:0] T781;
  wire[8:0] T782;
  wire T783;
  wire T784;
  reg [8:0] savedOffsets_19;
  wire[8:0] T927;
  wire[8:0] T785;
  wire[8:0] T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire T373;
  wire spillEndVal;
  wire T374;
  reg  spillEnd;
  wire T928;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire offsetUpdateVal_0;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire nextIterStartVal;
  wire T387;
  reg  nextIterStart;
  wire T929;
  wire T388;
  reg  offsetUpdate_0;
  wire T930;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire[31:0] T395;
  wire[4:0] T396;
  wire offsetUpdateVal_1;
  wire T397;
  wire T398;
  reg  offsetUpdate_1;
  wire T931;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire offsetUpdateVal_2;
  wire T405;
  wire T406;
  reg  offsetUpdate_2;
  wire T932;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire offsetUpdateVal_3;
  wire T411;
  wire T412;
  reg  offsetUpdate_3;
  wire T933;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire offsetUpdateVal_4;
  wire T421;
  wire T422;
  reg  offsetUpdate_4;
  wire T934;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire offsetUpdateVal_5;
  wire T427;
  wire T428;
  reg  offsetUpdate_5;
  wire T935;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire offsetUpdateVal_6;
  wire T435;
  wire T436;
  reg  offsetUpdate_6;
  wire T936;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire offsetUpdateVal_7;
  wire T441;
  wire T442;
  reg  offsetUpdate_7;
  wire T937;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire offsetUpdateVal_8;
  wire T453;
  wire T454;
  reg  offsetUpdate_8;
  wire T938;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire offsetUpdateVal_9;
  wire T459;
  wire T460;
  reg  offsetUpdate_9;
  wire T939;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire offsetUpdateVal_10;
  wire T467;
  wire T468;
  reg  offsetUpdate_10;
  wire T940;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire offsetUpdateVal_11;
  wire T473;
  wire T474;
  reg  offsetUpdate_11;
  wire T941;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire offsetUpdateVal_12;
  wire T483;
  wire T484;
  reg  offsetUpdate_12;
  wire T942;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire offsetUpdateVal_13;
  wire T489;
  wire T490;
  reg  offsetUpdate_13;
  wire T943;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire offsetUpdateVal_14;
  wire T497;
  wire T498;
  reg  offsetUpdate_14;
  wire T944;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire offsetUpdateVal_15;
  wire T503;
  wire T504;
  reg  offsetUpdate_15;
  wire T945;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire offsetUpdateVal_16;
  wire T515;
  wire T516;
  reg  offsetUpdate_16;
  wire T946;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire offsetUpdateVal_17;
  wire T521;
  wire T522;
  reg  offsetUpdate_17;
  wire T947;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire offsetUpdateVal_18;
  wire T529;
  wire T530;
  reg  offsetUpdate_18;
  wire T948;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire offsetUpdateVal_19;
  wire T535;
  wire T536;
  reg  offsetUpdate_19;
  wire T949;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire noCopyBaseAddrVal;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  reg  noCopyBaseAddr_0;
  wire T950;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire[31:0] T555;
  wire[4:0] T556;
  wire T557;
  wire T558;
  reg  noCopyBaseAddr_1;
  wire T951;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  reg  noCopyBaseAddr_2;
  wire T952;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  reg  noCopyBaseAddr_3;
  wire T953;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire T576;
  reg  noCopyBaseAddr_4;
  wire T954;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  reg  noCopyBaseAddr_5;
  wire T955;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  reg  noCopyBaseAddr_6;
  wire T956;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  reg  noCopyBaseAddr_7;
  wire T957;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  reg  noCopyBaseAddr_8;
  wire T958;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  reg  noCopyBaseAddr_9;
  wire T959;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  reg  noCopyBaseAddr_10;
  wire T960;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  reg  noCopyBaseAddr_11;
  wire T961;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  reg  noCopyBaseAddr_12;
  wire T962;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  reg  noCopyBaseAddr_13;
  wire T963;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  reg  noCopyBaseAddr_14;
  wire T964;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  reg  noCopyBaseAddr_15;
  wire T965;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  reg  noCopyBaseAddr_16;
  wire T966;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  reg  noCopyBaseAddr_17;
  wire T967;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  reg  noCopyBaseAddr_18;
  wire T968;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  reg  noCopyBaseAddr_19;
  wire T969;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[31:0] T668;
  wire[31:0] loopOffsetLkup;
  wire[31:0] T669;
  wire[31:0] T970;
  wire T670;
  wire T671;
  wire[31:0] T971;
  wire T792;
  wire T793;
  wire[31:0] T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire[31:0] T799;
  wire T800;
  wire T801;
  wire[31:0] baseAddrLkup;
  wire[31:0] T802;
  wire T803;
  wire T804;
  wire[63:0] T805;
  wire[63:0] T806;
  wire[63:0] T807;
  wire[63:0] T808;
  wire[63:0] T809;
  wire[63:0] T810;
  wire[63:0] T811;
  wire[63:0] T812;
  wire[63:0] T813;
  wire[63:0] T814;
  wire[63:0] T815;
  wire[63:0] T816;
  wire[63:0] T817;
  wire[63:0] T818;
  wire[63:0] T819;
  wire[63:0] T820;
  wire[63:0] T821;
  wire[63:0] T822;
  wire[63:0] T823;
  wire[4:0] T824;
  wire T825;
  wire[4:0] T826;
  wire T827;
  wire[8:0] T828;
  wire T829;
  wire[4:0] T830;
  wire T831;
  wire computeDone;
  wire T832;
  wire T833;
  wire T834;
  reg [2:0] compDoneCnt;
  wire[2:0] T972;
  wire[2:0] T835;
  wire[2:0] T836;
  wire[2:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire[63:0] T880;
  wire[31:0] baseAddrMem_io_outData;
  wire[42:0] storeSeqMem_io_outData;
  wire[31:0] loopOffsetMem_io_outData;
  wire[31:0] spillOffsetMem_io_outData;
  wire[8:0] storeSeqMemConfig_io_memAddr;
  wire[42:0] storeSeqMemConfig_io_memData;
  wire storeSeqMemConfig_io_memOutValid;
  wire storeSeqMemConfig_io_rst;
  wire[4:0] baseAddrMemConfig_io_memAddr;
  wire[31:0] baseAddrMemConfig_io_memData;
  wire baseAddrMemConfig_io_memOutValid;
  wire[4:0] loopOffsetMemConfig_io_memAddr;
  wire[31:0] loopOffsetMemConfig_io_memData;
  wire loopOffsetMemConfig_io_memOutValid;
  wire[4:0] spillOffsetMemConfig_io_memAddr;
  wire[31:0] spillOffsetMemConfig_io_memData;
  wire spillOffsetMemConfig_io_memOutValid;
  wire[63:0] storeReqFifo_io_deqData;
  wire storeReqFifo_io_enqRdy;
  wire storeReqFifo_io_deqValid;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    portSel_0 = {1{$random}};
    nextSeq = {2{$random}};
    nextSeqValid = {1{$random}};
    firstReqDone = {1{$random}};
    portSel_1 = {1{$random}};
    portSel_2 = {1{$random}};
    portSel_3 = {1{$random}};
    portSel_4 = {1{$random}};
    portSel_5 = {1{$random}};
    portSel_6 = {1{$random}};
    portSel_7 = {1{$random}};
    portSel_8 = {1{$random}};
    portSel_9 = {1{$random}};
    portSel_10 = {1{$random}};
    portSel_11 = {1{$random}};
    portSel_12 = {1{$random}};
    portSel_13 = {1{$random}};
    portSel_14 = {1{$random}};
    portSel_15 = {1{$random}};
    portSel_16 = {1{$random}};
    portSel_17 = {1{$random}};
    portSel_18 = {1{$random}};
    portSel_19 = {1{$random}};
    storeMemAddr = {1{$random}};
    savedOffsets_0 = {1{$random}};
    savedOffsets_1 = {1{$random}};
    savedOffsets_2 = {1{$random}};
    savedOffsets_3 = {1{$random}};
    savedOffsets_4 = {1{$random}};
    savedOffsets_5 = {1{$random}};
    savedOffsets_6 = {1{$random}};
    savedOffsets_7 = {1{$random}};
    savedOffsets_8 = {1{$random}};
    savedOffsets_9 = {1{$random}};
    savedOffsets_10 = {1{$random}};
    savedOffsets_11 = {1{$random}};
    savedOffsets_12 = {1{$random}};
    savedOffsets_13 = {1{$random}};
    savedOffsets_14 = {1{$random}};
    savedOffsets_15 = {1{$random}};
    savedOffsets_16 = {1{$random}};
    savedOffsets_17 = {1{$random}};
    savedOffsets_18 = {1{$random}};
    savedOffsets_19 = {1{$random}};
    spillEnd = {1{$random}};
    nextIterStart = {1{$random}};
    offsetUpdate_0 = {1{$random}};
    offsetUpdate_1 = {1{$random}};
    offsetUpdate_2 = {1{$random}};
    offsetUpdate_3 = {1{$random}};
    offsetUpdate_4 = {1{$random}};
    offsetUpdate_5 = {1{$random}};
    offsetUpdate_6 = {1{$random}};
    offsetUpdate_7 = {1{$random}};
    offsetUpdate_8 = {1{$random}};
    offsetUpdate_9 = {1{$random}};
    offsetUpdate_10 = {1{$random}};
    offsetUpdate_11 = {1{$random}};
    offsetUpdate_12 = {1{$random}};
    offsetUpdate_13 = {1{$random}};
    offsetUpdate_14 = {1{$random}};
    offsetUpdate_15 = {1{$random}};
    offsetUpdate_16 = {1{$random}};
    offsetUpdate_17 = {1{$random}};
    offsetUpdate_18 = {1{$random}};
    offsetUpdate_19 = {1{$random}};
    noCopyBaseAddr_0 = {1{$random}};
    noCopyBaseAddr_1 = {1{$random}};
    noCopyBaseAddr_2 = {1{$random}};
    noCopyBaseAddr_3 = {1{$random}};
    noCopyBaseAddr_4 = {1{$random}};
    noCopyBaseAddr_5 = {1{$random}};
    noCopyBaseAddr_6 = {1{$random}};
    noCopyBaseAddr_7 = {1{$random}};
    noCopyBaseAddr_8 = {1{$random}};
    noCopyBaseAddr_9 = {1{$random}};
    noCopyBaseAddr_10 = {1{$random}};
    noCopyBaseAddr_11 = {1{$random}};
    noCopyBaseAddr_12 = {1{$random}};
    noCopyBaseAddr_13 = {1{$random}};
    noCopyBaseAddr_14 = {1{$random}};
    noCopyBaseAddr_15 = {1{$random}};
    noCopyBaseAddr_16 = {1{$random}};
    noCopyBaseAddr_17 = {1{$random}};
    noCopyBaseAddr_18 = {1{$random}};
    noCopyBaseAddr_19 = {1{$random}};
    compDoneCnt = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = storeSeqMemConfig_io_rst ? 1'h1 : 1'h0;
  assign T1 = T231 ? 1'h0 : T2;
  assign T2 = T225 ? 1'h1 : T3;
  assign T3 = T224 ? 1'h0 : T4;
  assign T4 = T218 ? 1'h1 : T5;
  assign T5 = T217 ? 1'h0 : T6;
  assign T6 = T211 ? 1'h1 : T7;
  assign T7 = T210 ? 1'h0 : T8;
  assign T8 = T204 ? 1'h1 : T9;
  assign T9 = T203 ? 1'h0 : T10;
  assign T10 = T197 ? 1'h1 : T11;
  assign T11 = T196 ? 1'h0 : T12;
  assign T12 = T190 ? 1'h1 : T13;
  assign T13 = T189 ? 1'h0 : T14;
  assign T14 = T183 ? 1'h1 : T15;
  assign T15 = T182 ? 1'h0 : T16;
  assign T16 = T176 ? 1'h1 : T17;
  assign T17 = T175 ? 1'h0 : T18;
  assign T18 = T169 ? 1'h1 : T19;
  assign T19 = T168 ? 1'h0 : T20;
  assign T20 = T162 ? 1'h1 : T21;
  assign T21 = T161 ? 1'h0 : T22;
  assign T22 = T155 ? 1'h1 : T23;
  assign T23 = T154 ? 1'h0 : T24;
  assign T24 = T148 ? 1'h1 : T25;
  assign T25 = T147 ? 1'h0 : T26;
  assign T26 = T141 ? 1'h1 : T27;
  assign T27 = T140 ? 1'h0 : T28;
  assign T28 = T134 ? 1'h1 : T29;
  assign T29 = T133 ? 1'h0 : T30;
  assign T30 = T127 ? 1'h1 : T31;
  assign T31 = T126 ? 1'h0 : T32;
  assign T32 = T120 ? 1'h1 : T33;
  assign T33 = T119 ? 1'h0 : T34;
  assign T34 = T113 ? 1'h1 : T35;
  assign T35 = T112 ? 1'h0 : T36;
  assign T36 = T106 ? 1'h1 : T37;
  assign T37 = T105 ? 1'h0 : T38;
  assign T38 = T99 ? 1'h1 : T39;
  assign T39 = T40 ? 1'h1 : 1'h0;
  assign T40 = T41 & storeReqFifo_io_enqRdy;
  assign T41 = portSel_0 & io_fabOutToStoreValid_0;
  assign T881 = reset ? 1'h0 : T42;
  assign T42 = T40 ? 1'h0 : T43;
  assign T43 = T44 ? 1'h1 : portSel_0;
  assign T44 = T51 & T45;
  assign T45 = T46[1'h0:1'h0];
  assign T46 = 1'h1 << T47;
  assign T47 = portID;
  assign portID = T48;
  assign T48 = T51 ? T49 : 5'h0;
  assign T49 = nextSeq[6'h29:6'h25];
  assign T882 = reset ? 43'h0 : T50;
  assign T50 = io_seqMemAddrValid ? storeSeqMem_io_outData : nextSeq;
  assign T51 = T55 & nextSeqValid;
  assign T883 = reset ? 1'h0 : T52;
  assign T52 = T51 ? 1'h0 : T53;
  assign T53 = storeSeqMemConfig_io_rst ? 1'h0 : T54;
  assign T54 = io_seqMemAddrValid ? 1'h1 : nextSeqValid;
  assign T55 = getNextReq | T56;
  assign T56 = firstReqDone ^ 1'h1;
  assign T884 = reset ? 1'h0 : T57;
  assign T57 = T51 ? 1'h1 : T58;
  assign T58 = storeSeqMemConfig_io_rst ? 1'h0 : firstReqDone;
  assign getNextReq = T59;
  assign T59 = T231 ? 1'h0 : T60;
  assign T60 = T225 ? 1'h1 : T61;
  assign T61 = T224 ? 1'h0 : T62;
  assign T62 = T218 ? 1'h1 : T63;
  assign T63 = T217 ? 1'h0 : T64;
  assign T64 = T211 ? 1'h1 : T65;
  assign T65 = T210 ? 1'h0 : T66;
  assign T66 = T204 ? 1'h1 : T67;
  assign T67 = T203 ? 1'h0 : T68;
  assign T68 = T197 ? 1'h1 : T69;
  assign T69 = T196 ? 1'h0 : T70;
  assign T70 = T190 ? 1'h1 : T71;
  assign T71 = T189 ? 1'h0 : T72;
  assign T72 = T183 ? 1'h1 : T73;
  assign T73 = T182 ? 1'h0 : T74;
  assign T74 = T176 ? 1'h1 : T75;
  assign T75 = T175 ? 1'h0 : T76;
  assign T76 = T169 ? 1'h1 : T77;
  assign T77 = T168 ? 1'h0 : T78;
  assign T78 = T162 ? 1'h1 : T79;
  assign T79 = T161 ? 1'h0 : T80;
  assign T80 = T155 ? 1'h1 : T81;
  assign T81 = T154 ? 1'h0 : T82;
  assign T82 = T148 ? 1'h1 : T83;
  assign T83 = T147 ? 1'h0 : T84;
  assign T84 = T141 ? 1'h1 : T85;
  assign T85 = T140 ? 1'h0 : T86;
  assign T86 = T134 ? 1'h1 : T87;
  assign T87 = T133 ? 1'h0 : T88;
  assign T88 = T127 ? 1'h1 : T89;
  assign T89 = T126 ? 1'h0 : T90;
  assign T90 = T120 ? 1'h1 : T91;
  assign T91 = T119 ? 1'h0 : T92;
  assign T92 = T113 ? 1'h1 : T93;
  assign T93 = T112 ? 1'h0 : T94;
  assign T94 = T106 ? 1'h1 : T95;
  assign T95 = T105 ? 1'h0 : T96;
  assign T96 = T99 ? 1'h1 : T97;
  assign T97 = T98 ? 1'h0 : T40;
  assign T98 = T40 ^ 1'h1;
  assign T99 = T100 & storeReqFifo_io_enqRdy;
  assign T100 = portSel_1 & io_fabOutToStoreValid_1;
  assign T885 = reset ? 1'h0 : T101;
  assign T101 = T99 ? 1'h0 : T102;
  assign T102 = T103 ? 1'h1 : portSel_1;
  assign T103 = T51 & T104;
  assign T104 = T46[1'h1:1'h1];
  assign T105 = T99 ^ 1'h1;
  assign T106 = T107 & storeReqFifo_io_enqRdy;
  assign T107 = portSel_2 & io_fabOutToStoreValid_2;
  assign T886 = reset ? 1'h0 : T108;
  assign T108 = T106 ? 1'h0 : T109;
  assign T109 = T110 ? 1'h1 : portSel_2;
  assign T110 = T51 & T111;
  assign T111 = T46[2'h2:2'h2];
  assign T112 = T106 ^ 1'h1;
  assign T113 = T114 & storeReqFifo_io_enqRdy;
  assign T114 = portSel_3 & io_fabOutToStoreValid_3;
  assign T887 = reset ? 1'h0 : T115;
  assign T115 = T113 ? 1'h0 : T116;
  assign T116 = T117 ? 1'h1 : portSel_3;
  assign T117 = T51 & T118;
  assign T118 = T46[2'h3:2'h3];
  assign T119 = T113 ^ 1'h1;
  assign T120 = T121 & storeReqFifo_io_enqRdy;
  assign T121 = portSel_4 & io_fabOutToStoreValid_4;
  assign T888 = reset ? 1'h0 : T122;
  assign T122 = T120 ? 1'h0 : T123;
  assign T123 = T124 ? 1'h1 : portSel_4;
  assign T124 = T51 & T125;
  assign T125 = T46[3'h4:3'h4];
  assign T126 = T120 ^ 1'h1;
  assign T127 = T128 & storeReqFifo_io_enqRdy;
  assign T128 = portSel_5 & io_fabOutToStoreValid_5;
  assign T889 = reset ? 1'h0 : T129;
  assign T129 = T127 ? 1'h0 : T130;
  assign T130 = T131 ? 1'h1 : portSel_5;
  assign T131 = T51 & T132;
  assign T132 = T46[3'h5:3'h5];
  assign T133 = T127 ^ 1'h1;
  assign T134 = T135 & storeReqFifo_io_enqRdy;
  assign T135 = portSel_6 & io_fabOutToStoreValid_6;
  assign T890 = reset ? 1'h0 : T136;
  assign T136 = T134 ? 1'h0 : T137;
  assign T137 = T138 ? 1'h1 : portSel_6;
  assign T138 = T51 & T139;
  assign T139 = T46[3'h6:3'h6];
  assign T140 = T134 ^ 1'h1;
  assign T141 = T142 & storeReqFifo_io_enqRdy;
  assign T142 = portSel_7 & io_fabOutToStoreValid_7;
  assign T891 = reset ? 1'h0 : T143;
  assign T143 = T141 ? 1'h0 : T144;
  assign T144 = T145 ? 1'h1 : portSel_7;
  assign T145 = T51 & T146;
  assign T146 = T46[3'h7:3'h7];
  assign T147 = T141 ^ 1'h1;
  assign T148 = T149 & storeReqFifo_io_enqRdy;
  assign T149 = portSel_8 & io_fabOutToStoreValid_8;
  assign T892 = reset ? 1'h0 : T150;
  assign T150 = T148 ? 1'h0 : T151;
  assign T151 = T152 ? 1'h1 : portSel_8;
  assign T152 = T51 & T153;
  assign T153 = T46[4'h8:4'h8];
  assign T154 = T148 ^ 1'h1;
  assign T155 = T156 & storeReqFifo_io_enqRdy;
  assign T156 = portSel_9 & io_fabOutToStoreValid_9;
  assign T893 = reset ? 1'h0 : T157;
  assign T157 = T155 ? 1'h0 : T158;
  assign T158 = T159 ? 1'h1 : portSel_9;
  assign T159 = T51 & T160;
  assign T160 = T46[4'h9:4'h9];
  assign T161 = T155 ^ 1'h1;
  assign T162 = T163 & storeReqFifo_io_enqRdy;
  assign T163 = portSel_10 & io_fabOutToStoreValid_10;
  assign T894 = reset ? 1'h0 : T164;
  assign T164 = T162 ? 1'h0 : T165;
  assign T165 = T166 ? 1'h1 : portSel_10;
  assign T166 = T51 & T167;
  assign T167 = T46[4'ha:4'ha];
  assign T168 = T162 ^ 1'h1;
  assign T169 = T170 & storeReqFifo_io_enqRdy;
  assign T170 = portSel_11 & io_fabOutToStoreValid_11;
  assign T895 = reset ? 1'h0 : T171;
  assign T171 = T169 ? 1'h0 : T172;
  assign T172 = T173 ? 1'h1 : portSel_11;
  assign T173 = T51 & T174;
  assign T174 = T46[4'hb:4'hb];
  assign T175 = T169 ^ 1'h1;
  assign T176 = T177 & storeReqFifo_io_enqRdy;
  assign T177 = portSel_12 & io_fabOutToStoreValid_12;
  assign T896 = reset ? 1'h0 : T178;
  assign T178 = T176 ? 1'h0 : T179;
  assign T179 = T180 ? 1'h1 : portSel_12;
  assign T180 = T51 & T181;
  assign T181 = T46[4'hc:4'hc];
  assign T182 = T176 ^ 1'h1;
  assign T183 = T184 & storeReqFifo_io_enqRdy;
  assign T184 = portSel_13 & io_fabOutToStoreValid_13;
  assign T897 = reset ? 1'h0 : T185;
  assign T185 = T183 ? 1'h0 : T186;
  assign T186 = T187 ? 1'h1 : portSel_13;
  assign T187 = T51 & T188;
  assign T188 = T46[4'hd:4'hd];
  assign T189 = T183 ^ 1'h1;
  assign T190 = T191 & storeReqFifo_io_enqRdy;
  assign T191 = portSel_14 & io_fabOutToStoreValid_14;
  assign T898 = reset ? 1'h0 : T192;
  assign T192 = T190 ? 1'h0 : T193;
  assign T193 = T194 ? 1'h1 : portSel_14;
  assign T194 = T51 & T195;
  assign T195 = T46[4'he:4'he];
  assign T196 = T190 ^ 1'h1;
  assign T197 = T198 & storeReqFifo_io_enqRdy;
  assign T198 = portSel_15 & io_fabOutToStoreValid_15;
  assign T899 = reset ? 1'h0 : T199;
  assign T199 = T197 ? 1'h0 : T200;
  assign T200 = T201 ? 1'h1 : portSel_15;
  assign T201 = T51 & T202;
  assign T202 = T46[4'hf:4'hf];
  assign T203 = T197 ^ 1'h1;
  assign T204 = T205 & storeReqFifo_io_enqRdy;
  assign T205 = portSel_16 & io_fabOutToStoreValid_16;
  assign T900 = reset ? 1'h0 : T206;
  assign T206 = T204 ? 1'h0 : T207;
  assign T207 = T208 ? 1'h1 : portSel_16;
  assign T208 = T51 & T209;
  assign T209 = T46[5'h10:5'h10];
  assign T210 = T204 ^ 1'h1;
  assign T211 = T212 & storeReqFifo_io_enqRdy;
  assign T212 = portSel_17 & io_fabOutToStoreValid_17;
  assign T901 = reset ? 1'h0 : T213;
  assign T213 = T211 ? 1'h0 : T214;
  assign T214 = T215 ? 1'h1 : portSel_17;
  assign T215 = T51 & T216;
  assign T216 = T46[5'h11:5'h11];
  assign T217 = T211 ^ 1'h1;
  assign T218 = T219 & storeReqFifo_io_enqRdy;
  assign T219 = portSel_18 & io_fabOutToStoreValid_18;
  assign T902 = reset ? 1'h0 : T220;
  assign T220 = T218 ? 1'h0 : T221;
  assign T221 = T222 ? 1'h1 : portSel_18;
  assign T222 = T51 & T223;
  assign T223 = T46[5'h12:5'h12];
  assign T224 = T218 ^ 1'h1;
  assign T225 = T226 & storeReqFifo_io_enqRdy;
  assign T226 = portSel_19 & io_fabOutToStoreValid_19;
  assign T903 = reset ? 1'h0 : T227;
  assign T227 = T225 ? 1'h0 : T228;
  assign T228 = T229 ? 1'h1 : portSel_19;
  assign T229 = T51 & T230;
  assign T230 = T46[5'h13:5'h13];
  assign T231 = T225 ^ 1'h1;
  assign T232 = io_storeMemRdy ? io_storeMemRdy : io_storeMemRdy;
  assign T233 = T231 ? 64'h0 : T234;
  assign T234 = T225 ? T823 : T235;
  assign T235 = T224 ? 64'h0 : T236;
  assign T236 = T218 ? T822 : T237;
  assign T237 = T217 ? 64'h0 : T238;
  assign T238 = T211 ? T821 : T239;
  assign T239 = T210 ? 64'h0 : T240;
  assign T240 = T204 ? T820 : T241;
  assign T241 = T203 ? 64'h0 : T242;
  assign T242 = T197 ? T819 : T243;
  assign T243 = T196 ? 64'h0 : T244;
  assign T244 = T190 ? T818 : T245;
  assign T245 = T189 ? 64'h0 : T246;
  assign T246 = T183 ? T817 : T247;
  assign T247 = T182 ? 64'h0 : T248;
  assign T248 = T176 ? T816 : T249;
  assign T249 = T175 ? 64'h0 : T250;
  assign T250 = T169 ? T815 : T251;
  assign T251 = T168 ? 64'h0 : T252;
  assign T252 = T162 ? T814 : T253;
  assign T253 = T161 ? 64'h0 : T254;
  assign T254 = T155 ? T813 : T255;
  assign T255 = T154 ? 64'h0 : T256;
  assign T256 = T148 ? T812 : T257;
  assign T257 = T147 ? 64'h0 : T258;
  assign T258 = T141 ? T811 : T259;
  assign T259 = T140 ? 64'h0 : T260;
  assign T260 = T134 ? T810 : T261;
  assign T261 = T133 ? 64'h0 : T262;
  assign T262 = T127 ? T809 : T263;
  assign T263 = T126 ? 64'h0 : T264;
  assign T264 = T120 ? T808 : T265;
  assign T265 = T119 ? 64'h0 : T266;
  assign T266 = T113 ? T807 : T267;
  assign T267 = T112 ? 64'h0 : T268;
  assign T268 = T106 ? T806 : T269;
  assign T269 = T105 ? 64'h0 : T270;
  assign T270 = T99 ? T805 : T271;
  assign T271 = T40 ? T272 : 64'h0;
  assign T272 = {storeReqAddr, storeReqData};
  assign storeReqData = T273;
  assign T273 = T231 ? 32'h0 : T274;
  assign T274 = T225 ? io_fabOutToStore_19 : T275;
  assign T275 = T224 ? 32'h0 : T276;
  assign T276 = T218 ? io_fabOutToStore_18 : T277;
  assign T277 = T217 ? 32'h0 : T278;
  assign T278 = T211 ? io_fabOutToStore_17 : T279;
  assign T279 = T210 ? 32'h0 : T280;
  assign T280 = T204 ? io_fabOutToStore_16 : T281;
  assign T281 = T203 ? 32'h0 : T282;
  assign T282 = T197 ? io_fabOutToStore_15 : T283;
  assign T283 = T196 ? 32'h0 : T284;
  assign T284 = T190 ? io_fabOutToStore_14 : T285;
  assign T285 = T189 ? 32'h0 : T286;
  assign T286 = T183 ? io_fabOutToStore_13 : T287;
  assign T287 = T182 ? 32'h0 : T288;
  assign T288 = T176 ? io_fabOutToStore_12 : T289;
  assign T289 = T175 ? 32'h0 : T290;
  assign T290 = T169 ? io_fabOutToStore_11 : T291;
  assign T291 = T168 ? 32'h0 : T292;
  assign T292 = T162 ? io_fabOutToStore_10 : T293;
  assign T293 = T161 ? 32'h0 : T294;
  assign T294 = T155 ? io_fabOutToStore_9 : T295;
  assign T295 = T154 ? 32'h0 : T296;
  assign T296 = T148 ? io_fabOutToStore_8 : T297;
  assign T297 = T147 ? 32'h0 : T298;
  assign T298 = T141 ? io_fabOutToStore_7 : T299;
  assign T299 = T140 ? 32'h0 : T300;
  assign T300 = T134 ? io_fabOutToStore_6 : T301;
  assign T301 = T133 ? 32'h0 : T302;
  assign T302 = T127 ? io_fabOutToStore_5 : T303;
  assign T303 = T126 ? 32'h0 : T304;
  assign T304 = T120 ? io_fabOutToStore_4 : T305;
  assign T305 = T119 ? 32'h0 : T306;
  assign T306 = T113 ? io_fabOutToStore_3 : T307;
  assign T307 = T112 ? 32'h0 : T308;
  assign T308 = T106 ? io_fabOutToStore_2 : T309;
  assign T309 = T105 ? 32'h0 : T310;
  assign T310 = T99 ? io_fabOutToStore_1 : T311;
  assign T311 = T98 ? 32'h0 : T312;
  assign T312 = T40 ? io_fabOutToStore_0 : 32'h0;
  assign storeReqAddr = T313;
  assign T313 = T231 ? 32'h0 : T314;
  assign T314 = T225 ? storeMemAddr : T315;
  assign T315 = T224 ? 32'h0 : T316;
  assign T316 = T218 ? storeMemAddr : T317;
  assign T317 = T217 ? 32'h0 : T318;
  assign T318 = T211 ? storeMemAddr : T319;
  assign T319 = T210 ? 32'h0 : T320;
  assign T320 = T204 ? storeMemAddr : T321;
  assign T321 = T203 ? 32'h0 : T322;
  assign T322 = T197 ? storeMemAddr : T323;
  assign T323 = T196 ? 32'h0 : T324;
  assign T324 = T190 ? storeMemAddr : T325;
  assign T325 = T189 ? 32'h0 : T326;
  assign T326 = T183 ? storeMemAddr : T327;
  assign T327 = T182 ? 32'h0 : T328;
  assign T328 = T176 ? storeMemAddr : T329;
  assign T329 = T175 ? 32'h0 : T330;
  assign T330 = T169 ? storeMemAddr : T331;
  assign T331 = T168 ? 32'h0 : T332;
  assign T332 = T162 ? storeMemAddr : T333;
  assign T333 = T161 ? 32'h0 : T334;
  assign T334 = T155 ? storeMemAddr : T335;
  assign T335 = T154 ? 32'h0 : T336;
  assign T336 = T148 ? storeMemAddr : T337;
  assign T337 = T147 ? 32'h0 : T338;
  assign T338 = T141 ? storeMemAddr : T339;
  assign T339 = T140 ? 32'h0 : T340;
  assign T340 = T134 ? storeMemAddr : T341;
  assign T341 = T133 ? 32'h0 : T342;
  assign T342 = T127 ? storeMemAddr : T343;
  assign T343 = T126 ? 32'h0 : T344;
  assign T344 = T120 ? storeMemAddr : T345;
  assign T345 = T119 ? 32'h0 : T346;
  assign T346 = T113 ? storeMemAddr : T347;
  assign T347 = T112 ? 32'h0 : T348;
  assign T348 = T106 ? storeMemAddr : T349;
  assign T349 = T105 ? 32'h0 : T350;
  assign T350 = T99 ? storeMemAddr : T351;
  assign T351 = T98 ? 32'h0 : T352;
  assign T352 = T40 ? storeMemAddr : 32'h0;
  assign T904 = reset ? 32'h0 : T353;
  assign T353 = T51 ? T354 : storeMemAddr;
  assign T354 = T905 + offsetAddr;
  assign offsetAddr = T355;
  assign T355 = T51 ? T356 : 32'h0;
  assign T356 = nextSeq[6'h24:3'h5];
  assign T905 = {31'h0, T357};
  assign T357 = T364 & T358;
  assign T358 = T359 - 1'h1;
  assign T359 = 1'h1 << T360;
  assign T360 = T361 + 5'h1;
  assign T361 = addrLkupIndex - addrLkupIndex;
  assign addrLkupIndex = T362;
  assign T362 = T51 ? T363 : 5'h0;
  assign T363 = nextSeq[3'h4:1'h0];
  assign T364 = savedOffsetsVal >> addrLkupIndex;
  assign savedOffsetsVal = T906;
  assign T906 = T365[4'h8:1'h0];
  assign T365 = T803 ? baseAddrLkup : T366;
  assign T366 = T800 ? T799 : T367;
  assign T367 = T795 ? T794 : T368;
  assign T368 = T792 ? T971 : T369;
  assign T369 = T670 ? T668 : T370;
  assign T370 = T373 ? T371 : 32'h0;
  assign T371 = T907 - spillLkup;
  assign spillLkup = T372;
  assign T372 = T51 ? spillOffsetMem_io_outData : 32'h0;
  assign T907 = {23'h0, T672};
  assign T672 = T791 ? T769 : T673;
  assign T673 = T768 ? T722 : T674;
  assign T674 = T721 ? T699 : T675;
  assign T675 = T698 ? T688 : T676;
  assign T676 = T687 ? savedOffsets_1 : savedOffsets_0;
  assign T908 = reset ? 9'h0 : T677;
  assign T677 = T679 ? savedOffsetsVal : T678;
  assign T678 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_0;
  assign T679 = T51 & T680;
  assign T680 = T681[1'h0:1'h0];
  assign T681 = 1'h1 << T682;
  assign T682 = addrLkupIndex;
  assign T909 = reset ? 9'h0 : T683;
  assign T683 = T685 ? savedOffsetsVal : T684;
  assign T684 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_1;
  assign T685 = T51 & T686;
  assign T686 = T681[1'h1:1'h1];
  assign T687 = T682[1'h0:1'h0];
  assign T688 = T697 ? savedOffsets_3 : savedOffsets_2;
  assign T910 = reset ? 9'h0 : T689;
  assign T689 = T691 ? savedOffsetsVal : T690;
  assign T690 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_2;
  assign T691 = T51 & T692;
  assign T692 = T681[2'h2:2'h2];
  assign T911 = reset ? 9'h0 : T693;
  assign T693 = T695 ? savedOffsetsVal : T694;
  assign T694 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_3;
  assign T695 = T51 & T696;
  assign T696 = T681[2'h3:2'h3];
  assign T697 = T682[1'h0:1'h0];
  assign T698 = T682[1'h1:1'h1];
  assign T699 = T720 ? T710 : T700;
  assign T700 = T709 ? savedOffsets_5 : savedOffsets_4;
  assign T912 = reset ? 9'h0 : T701;
  assign T701 = T703 ? savedOffsetsVal : T702;
  assign T702 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_4;
  assign T703 = T51 & T704;
  assign T704 = T681[3'h4:3'h4];
  assign T913 = reset ? 9'h0 : T705;
  assign T705 = T707 ? savedOffsetsVal : T706;
  assign T706 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_5;
  assign T707 = T51 & T708;
  assign T708 = T681[3'h5:3'h5];
  assign T709 = T682[1'h0:1'h0];
  assign T710 = T719 ? savedOffsets_7 : savedOffsets_6;
  assign T914 = reset ? 9'h0 : T711;
  assign T711 = T713 ? savedOffsetsVal : T712;
  assign T712 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_6;
  assign T713 = T51 & T714;
  assign T714 = T681[3'h6:3'h6];
  assign T915 = reset ? 9'h0 : T715;
  assign T715 = T717 ? savedOffsetsVal : T716;
  assign T716 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_7;
  assign T717 = T51 & T718;
  assign T718 = T681[3'h7:3'h7];
  assign T719 = T682[1'h0:1'h0];
  assign T720 = T682[1'h1:1'h1];
  assign T721 = T682[2'h2:2'h2];
  assign T722 = T767 ? T745 : T723;
  assign T723 = T744 ? T734 : T724;
  assign T724 = T733 ? savedOffsets_9 : savedOffsets_8;
  assign T916 = reset ? 9'h0 : T725;
  assign T725 = T727 ? savedOffsetsVal : T726;
  assign T726 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_8;
  assign T727 = T51 & T728;
  assign T728 = T681[4'h8:4'h8];
  assign T917 = reset ? 9'h0 : T729;
  assign T729 = T731 ? savedOffsetsVal : T730;
  assign T730 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_9;
  assign T731 = T51 & T732;
  assign T732 = T681[4'h9:4'h9];
  assign T733 = T682[1'h0:1'h0];
  assign T734 = T743 ? savedOffsets_11 : savedOffsets_10;
  assign T918 = reset ? 9'h0 : T735;
  assign T735 = T737 ? savedOffsetsVal : T736;
  assign T736 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_10;
  assign T737 = T51 & T738;
  assign T738 = T681[4'ha:4'ha];
  assign T919 = reset ? 9'h0 : T739;
  assign T739 = T741 ? savedOffsetsVal : T740;
  assign T740 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_11;
  assign T741 = T51 & T742;
  assign T742 = T681[4'hb:4'hb];
  assign T743 = T682[1'h0:1'h0];
  assign T744 = T682[1'h1:1'h1];
  assign T745 = T766 ? T756 : T746;
  assign T746 = T755 ? savedOffsets_13 : savedOffsets_12;
  assign T920 = reset ? 9'h0 : T747;
  assign T747 = T749 ? savedOffsetsVal : T748;
  assign T748 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_12;
  assign T749 = T51 & T750;
  assign T750 = T681[4'hc:4'hc];
  assign T921 = reset ? 9'h0 : T751;
  assign T751 = T753 ? savedOffsetsVal : T752;
  assign T752 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_13;
  assign T753 = T51 & T754;
  assign T754 = T681[4'hd:4'hd];
  assign T755 = T682[1'h0:1'h0];
  assign T756 = T765 ? savedOffsets_15 : savedOffsets_14;
  assign T922 = reset ? 9'h0 : T757;
  assign T757 = T759 ? savedOffsetsVal : T758;
  assign T758 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_14;
  assign T759 = T51 & T760;
  assign T760 = T681[4'he:4'he];
  assign T923 = reset ? 9'h0 : T761;
  assign T761 = T763 ? savedOffsetsVal : T762;
  assign T762 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_15;
  assign T763 = T51 & T764;
  assign T764 = T681[4'hf:4'hf];
  assign T765 = T682[1'h0:1'h0];
  assign T766 = T682[1'h1:1'h1];
  assign T767 = T682[2'h2:2'h2];
  assign T768 = T682[2'h3:2'h3];
  assign T769 = T790 ? T780 : T770;
  assign T770 = T779 ? savedOffsets_17 : savedOffsets_16;
  assign T924 = reset ? 9'h0 : T771;
  assign T771 = T773 ? savedOffsetsVal : T772;
  assign T772 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_16;
  assign T773 = T51 & T774;
  assign T774 = T681[5'h10:5'h10];
  assign T925 = reset ? 9'h0 : T775;
  assign T775 = T777 ? savedOffsetsVal : T776;
  assign T776 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_17;
  assign T777 = T51 & T778;
  assign T778 = T681[5'h11:5'h11];
  assign T779 = T682[1'h0:1'h0];
  assign T780 = T789 ? savedOffsets_19 : savedOffsets_18;
  assign T926 = reset ? 9'h0 : T781;
  assign T781 = T783 ? savedOffsetsVal : T782;
  assign T782 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_18;
  assign T783 = T51 & T784;
  assign T784 = T681[5'h12:5'h12];
  assign T927 = reset ? 9'h0 : T785;
  assign T785 = T787 ? savedOffsetsVal : T786;
  assign T786 = storeSeqMemConfig_io_rst ? 9'h0 : savedOffsets_19;
  assign T787 = T51 & T788;
  assign T788 = T681[5'h13:5'h13];
  assign T789 = T682[1'h0:1'h0];
  assign T790 = T682[1'h1:1'h1];
  assign T791 = T682[3'h4:3'h4];
  assign T373 = T377 & spillEndVal;
  assign spillEndVal = T374;
  assign T374 = T51 ? spillEnd : 1'h0;
  assign T928 = reset ? 1'h0 : T375;
  assign T375 = storeSeqMemConfig_io_rst ? 1'h0 : T376;
  assign T376 = io_seqMemAddrValid ? io_spillEnd : spillEnd;
  assign T377 = T544 & T378;
  assign T378 = T543 ? T513 : T379;
  assign T379 = T512 ? T450 : T380;
  assign T380 = T449 ? T419 : T381;
  assign T381 = T418 ? T404 : T382;
  assign T382 = T403 ? offsetUpdateVal_1 : offsetUpdateVal_0;
  assign offsetUpdateVal_0 = T383;
  assign T383 = T393 ? 1'h0 : T384;
  assign T384 = T391 ? offsetUpdate_0 : T385;
  assign T385 = T51 & T386;
  assign T386 = spillEndVal | nextIterStartVal;
  assign nextIterStartVal = T387;
  assign T387 = T51 ? nextIterStart : 1'h0;
  assign T929 = reset ? 1'h0 : T388;
  assign T388 = io_seqMemAddrValid ? io_nextIterStart : nextIterStart;
  assign T930 = reset ? 1'h0 : T389;
  assign T389 = T51 ? offsetUpdateVal_0 : T390;
  assign T390 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_0;
  assign T391 = T51 & T392;
  assign T392 = T386 ^ 1'h1;
  assign T393 = T51 & T394;
  assign T394 = T395[1'h0:1'h0];
  assign T395 = 1'h1 << T396;
  assign T396 = addrLkupIndex;
  assign offsetUpdateVal_1 = T397;
  assign T397 = T401 ? 1'h0 : T398;
  assign T398 = T391 ? offsetUpdate_1 : T385;
  assign T931 = reset ? 1'h0 : T399;
  assign T399 = T51 ? offsetUpdateVal_1 : T400;
  assign T400 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_1;
  assign T401 = T51 & T402;
  assign T402 = T395[1'h1:1'h1];
  assign T403 = T396[1'h0:1'h0];
  assign T404 = T417 ? offsetUpdateVal_3 : offsetUpdateVal_2;
  assign offsetUpdateVal_2 = T405;
  assign T405 = T409 ? 1'h0 : T406;
  assign T406 = T391 ? offsetUpdate_2 : T385;
  assign T932 = reset ? 1'h0 : T407;
  assign T407 = T51 ? offsetUpdateVal_2 : T408;
  assign T408 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_2;
  assign T409 = T51 & T410;
  assign T410 = T395[2'h2:2'h2];
  assign offsetUpdateVal_3 = T411;
  assign T411 = T415 ? 1'h0 : T412;
  assign T412 = T391 ? offsetUpdate_3 : T385;
  assign T933 = reset ? 1'h0 : T413;
  assign T413 = T51 ? offsetUpdateVal_3 : T414;
  assign T414 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_3;
  assign T415 = T51 & T416;
  assign T416 = T395[2'h3:2'h3];
  assign T417 = T396[1'h0:1'h0];
  assign T418 = T396[1'h1:1'h1];
  assign T419 = T448 ? T434 : T420;
  assign T420 = T433 ? offsetUpdateVal_5 : offsetUpdateVal_4;
  assign offsetUpdateVal_4 = T421;
  assign T421 = T425 ? 1'h0 : T422;
  assign T422 = T391 ? offsetUpdate_4 : T385;
  assign T934 = reset ? 1'h0 : T423;
  assign T423 = T51 ? offsetUpdateVal_4 : T424;
  assign T424 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_4;
  assign T425 = T51 & T426;
  assign T426 = T395[3'h4:3'h4];
  assign offsetUpdateVal_5 = T427;
  assign T427 = T431 ? 1'h0 : T428;
  assign T428 = T391 ? offsetUpdate_5 : T385;
  assign T935 = reset ? 1'h0 : T429;
  assign T429 = T51 ? offsetUpdateVal_5 : T430;
  assign T430 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_5;
  assign T431 = T51 & T432;
  assign T432 = T395[3'h5:3'h5];
  assign T433 = T396[1'h0:1'h0];
  assign T434 = T447 ? offsetUpdateVal_7 : offsetUpdateVal_6;
  assign offsetUpdateVal_6 = T435;
  assign T435 = T439 ? 1'h0 : T436;
  assign T436 = T391 ? offsetUpdate_6 : T385;
  assign T936 = reset ? 1'h0 : T437;
  assign T437 = T51 ? offsetUpdateVal_6 : T438;
  assign T438 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_6;
  assign T439 = T51 & T440;
  assign T440 = T395[3'h6:3'h6];
  assign offsetUpdateVal_7 = T441;
  assign T441 = T445 ? 1'h0 : T442;
  assign T442 = T391 ? offsetUpdate_7 : T385;
  assign T937 = reset ? 1'h0 : T443;
  assign T443 = T51 ? offsetUpdateVal_7 : T444;
  assign T444 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_7;
  assign T445 = T51 & T446;
  assign T446 = T395[3'h7:3'h7];
  assign T447 = T396[1'h0:1'h0];
  assign T448 = T396[1'h1:1'h1];
  assign T449 = T396[2'h2:2'h2];
  assign T450 = T511 ? T481 : T451;
  assign T451 = T480 ? T466 : T452;
  assign T452 = T465 ? offsetUpdateVal_9 : offsetUpdateVal_8;
  assign offsetUpdateVal_8 = T453;
  assign T453 = T457 ? 1'h0 : T454;
  assign T454 = T391 ? offsetUpdate_8 : T385;
  assign T938 = reset ? 1'h0 : T455;
  assign T455 = T51 ? offsetUpdateVal_8 : T456;
  assign T456 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_8;
  assign T457 = T51 & T458;
  assign T458 = T395[4'h8:4'h8];
  assign offsetUpdateVal_9 = T459;
  assign T459 = T463 ? 1'h0 : T460;
  assign T460 = T391 ? offsetUpdate_9 : T385;
  assign T939 = reset ? 1'h0 : T461;
  assign T461 = T51 ? offsetUpdateVal_9 : T462;
  assign T462 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_9;
  assign T463 = T51 & T464;
  assign T464 = T395[4'h9:4'h9];
  assign T465 = T396[1'h0:1'h0];
  assign T466 = T479 ? offsetUpdateVal_11 : offsetUpdateVal_10;
  assign offsetUpdateVal_10 = T467;
  assign T467 = T471 ? 1'h0 : T468;
  assign T468 = T391 ? offsetUpdate_10 : T385;
  assign T940 = reset ? 1'h0 : T469;
  assign T469 = T51 ? offsetUpdateVal_10 : T470;
  assign T470 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_10;
  assign T471 = T51 & T472;
  assign T472 = T395[4'ha:4'ha];
  assign offsetUpdateVal_11 = T473;
  assign T473 = T477 ? 1'h0 : T474;
  assign T474 = T391 ? offsetUpdate_11 : T385;
  assign T941 = reset ? 1'h0 : T475;
  assign T475 = T51 ? offsetUpdateVal_11 : T476;
  assign T476 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_11;
  assign T477 = T51 & T478;
  assign T478 = T395[4'hb:4'hb];
  assign T479 = T396[1'h0:1'h0];
  assign T480 = T396[1'h1:1'h1];
  assign T481 = T510 ? T496 : T482;
  assign T482 = T495 ? offsetUpdateVal_13 : offsetUpdateVal_12;
  assign offsetUpdateVal_12 = T483;
  assign T483 = T487 ? 1'h0 : T484;
  assign T484 = T391 ? offsetUpdate_12 : T385;
  assign T942 = reset ? 1'h0 : T485;
  assign T485 = T51 ? offsetUpdateVal_12 : T486;
  assign T486 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_12;
  assign T487 = T51 & T488;
  assign T488 = T395[4'hc:4'hc];
  assign offsetUpdateVal_13 = T489;
  assign T489 = T493 ? 1'h0 : T490;
  assign T490 = T391 ? offsetUpdate_13 : T385;
  assign T943 = reset ? 1'h0 : T491;
  assign T491 = T51 ? offsetUpdateVal_13 : T492;
  assign T492 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_13;
  assign T493 = T51 & T494;
  assign T494 = T395[4'hd:4'hd];
  assign T495 = T396[1'h0:1'h0];
  assign T496 = T509 ? offsetUpdateVal_15 : offsetUpdateVal_14;
  assign offsetUpdateVal_14 = T497;
  assign T497 = T501 ? 1'h0 : T498;
  assign T498 = T391 ? offsetUpdate_14 : T385;
  assign T944 = reset ? 1'h0 : T499;
  assign T499 = T51 ? offsetUpdateVal_14 : T500;
  assign T500 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_14;
  assign T501 = T51 & T502;
  assign T502 = T395[4'he:4'he];
  assign offsetUpdateVal_15 = T503;
  assign T503 = T507 ? 1'h0 : T504;
  assign T504 = T391 ? offsetUpdate_15 : T385;
  assign T945 = reset ? 1'h0 : T505;
  assign T505 = T51 ? offsetUpdateVal_15 : T506;
  assign T506 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_15;
  assign T507 = T51 & T508;
  assign T508 = T395[4'hf:4'hf];
  assign T509 = T396[1'h0:1'h0];
  assign T510 = T396[1'h1:1'h1];
  assign T511 = T396[2'h2:2'h2];
  assign T512 = T396[2'h3:2'h3];
  assign T513 = T542 ? T528 : T514;
  assign T514 = T527 ? offsetUpdateVal_17 : offsetUpdateVal_16;
  assign offsetUpdateVal_16 = T515;
  assign T515 = T519 ? 1'h0 : T516;
  assign T516 = T391 ? offsetUpdate_16 : T385;
  assign T946 = reset ? 1'h0 : T517;
  assign T517 = T51 ? offsetUpdateVal_16 : T518;
  assign T518 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_16;
  assign T519 = T51 & T520;
  assign T520 = T395[5'h10:5'h10];
  assign offsetUpdateVal_17 = T521;
  assign T521 = T525 ? 1'h0 : T522;
  assign T522 = T391 ? offsetUpdate_17 : T385;
  assign T947 = reset ? 1'h0 : T523;
  assign T523 = T51 ? offsetUpdateVal_17 : T524;
  assign T524 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_17;
  assign T525 = T51 & T526;
  assign T526 = T395[5'h11:5'h11];
  assign T527 = T396[1'h0:1'h0];
  assign T528 = T541 ? offsetUpdateVal_19 : offsetUpdateVal_18;
  assign offsetUpdateVal_18 = T529;
  assign T529 = T533 ? 1'h0 : T530;
  assign T530 = T391 ? offsetUpdate_18 : T385;
  assign T948 = reset ? 1'h0 : T531;
  assign T531 = T51 ? offsetUpdateVal_18 : T532;
  assign T532 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_18;
  assign T533 = T51 & T534;
  assign T534 = T395[5'h12:5'h12];
  assign offsetUpdateVal_19 = T535;
  assign T535 = T539 ? 1'h0 : T536;
  assign T536 = T391 ? offsetUpdate_19 : T385;
  assign T949 = reset ? 1'h0 : T537;
  assign T537 = T51 ? offsetUpdateVal_19 : T538;
  assign T538 = storeSeqMemConfig_io_rst ? 1'h0 : offsetUpdate_19;
  assign T539 = T51 & T540;
  assign T540 = T395[5'h13:5'h13];
  assign T541 = T396[1'h0:1'h0];
  assign T542 = T396[1'h1:1'h1];
  assign T543 = T396[3'h4:3'h4];
  assign T544 = T51 & noCopyBaseAddrVal;
  assign noCopyBaseAddrVal = T545;
  assign T545 = T51 ? T546 : 1'h0;
  assign T546 = T667 ? T645 : T547;
  assign T547 = T644 ? T598 : T548;
  assign T548 = T597 ? T575 : T549;
  assign T549 = T574 ? T564 : T550;
  assign T550 = T563 ? noCopyBaseAddr_1 : noCopyBaseAddr_0;
  assign T950 = reset ? 1'h0 : T551;
  assign T551 = T553 ? 1'h1 : T552;
  assign T552 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_0;
  assign T553 = T557 & T554;
  assign T554 = T555[1'h0:1'h0];
  assign T555 = 1'h1 << T556;
  assign T556 = addrLkupIndex;
  assign T557 = T51 & T558;
  assign T558 = noCopyBaseAddrVal ^ 1'h1;
  assign T951 = reset ? 1'h0 : T559;
  assign T559 = T561 ? 1'h1 : T560;
  assign T560 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_1;
  assign T561 = T557 & T562;
  assign T562 = T555[1'h1:1'h1];
  assign T563 = T556[1'h0:1'h0];
  assign T564 = T573 ? noCopyBaseAddr_3 : noCopyBaseAddr_2;
  assign T952 = reset ? 1'h0 : T565;
  assign T565 = T567 ? 1'h1 : T566;
  assign T566 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_2;
  assign T567 = T557 & T568;
  assign T568 = T555[2'h2:2'h2];
  assign T953 = reset ? 1'h0 : T569;
  assign T569 = T571 ? 1'h1 : T570;
  assign T570 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_3;
  assign T571 = T557 & T572;
  assign T572 = T555[2'h3:2'h3];
  assign T573 = T556[1'h0:1'h0];
  assign T574 = T556[1'h1:1'h1];
  assign T575 = T596 ? T586 : T576;
  assign T576 = T585 ? noCopyBaseAddr_5 : noCopyBaseAddr_4;
  assign T954 = reset ? 1'h0 : T577;
  assign T577 = T579 ? 1'h1 : T578;
  assign T578 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_4;
  assign T579 = T557 & T580;
  assign T580 = T555[3'h4:3'h4];
  assign T955 = reset ? 1'h0 : T581;
  assign T581 = T583 ? 1'h1 : T582;
  assign T582 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_5;
  assign T583 = T557 & T584;
  assign T584 = T555[3'h5:3'h5];
  assign T585 = T556[1'h0:1'h0];
  assign T586 = T595 ? noCopyBaseAddr_7 : noCopyBaseAddr_6;
  assign T956 = reset ? 1'h0 : T587;
  assign T587 = T589 ? 1'h1 : T588;
  assign T588 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_6;
  assign T589 = T557 & T590;
  assign T590 = T555[3'h6:3'h6];
  assign T957 = reset ? 1'h0 : T591;
  assign T591 = T593 ? 1'h1 : T592;
  assign T592 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_7;
  assign T593 = T557 & T594;
  assign T594 = T555[3'h7:3'h7];
  assign T595 = T556[1'h0:1'h0];
  assign T596 = T556[1'h1:1'h1];
  assign T597 = T556[2'h2:2'h2];
  assign T598 = T643 ? T621 : T599;
  assign T599 = T620 ? T610 : T600;
  assign T600 = T609 ? noCopyBaseAddr_9 : noCopyBaseAddr_8;
  assign T958 = reset ? 1'h0 : T601;
  assign T601 = T603 ? 1'h1 : T602;
  assign T602 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_8;
  assign T603 = T557 & T604;
  assign T604 = T555[4'h8:4'h8];
  assign T959 = reset ? 1'h0 : T605;
  assign T605 = T607 ? 1'h1 : T606;
  assign T606 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_9;
  assign T607 = T557 & T608;
  assign T608 = T555[4'h9:4'h9];
  assign T609 = T556[1'h0:1'h0];
  assign T610 = T619 ? noCopyBaseAddr_11 : noCopyBaseAddr_10;
  assign T960 = reset ? 1'h0 : T611;
  assign T611 = T613 ? 1'h1 : T612;
  assign T612 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_10;
  assign T613 = T557 & T614;
  assign T614 = T555[4'ha:4'ha];
  assign T961 = reset ? 1'h0 : T615;
  assign T615 = T617 ? 1'h1 : T616;
  assign T616 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_11;
  assign T617 = T557 & T618;
  assign T618 = T555[4'hb:4'hb];
  assign T619 = T556[1'h0:1'h0];
  assign T620 = T556[1'h1:1'h1];
  assign T621 = T642 ? T632 : T622;
  assign T622 = T631 ? noCopyBaseAddr_13 : noCopyBaseAddr_12;
  assign T962 = reset ? 1'h0 : T623;
  assign T623 = T625 ? 1'h1 : T624;
  assign T624 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_12;
  assign T625 = T557 & T626;
  assign T626 = T555[4'hc:4'hc];
  assign T963 = reset ? 1'h0 : T627;
  assign T627 = T629 ? 1'h1 : T628;
  assign T628 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_13;
  assign T629 = T557 & T630;
  assign T630 = T555[4'hd:4'hd];
  assign T631 = T556[1'h0:1'h0];
  assign T632 = T641 ? noCopyBaseAddr_15 : noCopyBaseAddr_14;
  assign T964 = reset ? 1'h0 : T633;
  assign T633 = T635 ? 1'h1 : T634;
  assign T634 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_14;
  assign T635 = T557 & T636;
  assign T636 = T555[4'he:4'he];
  assign T965 = reset ? 1'h0 : T637;
  assign T637 = T639 ? 1'h1 : T638;
  assign T638 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_15;
  assign T639 = T557 & T640;
  assign T640 = T555[4'hf:4'hf];
  assign T641 = T556[1'h0:1'h0];
  assign T642 = T556[1'h1:1'h1];
  assign T643 = T556[2'h2:2'h2];
  assign T644 = T556[2'h3:2'h3];
  assign T645 = T666 ? T656 : T646;
  assign T646 = T655 ? noCopyBaseAddr_17 : noCopyBaseAddr_16;
  assign T966 = reset ? 1'h0 : T647;
  assign T647 = T649 ? 1'h1 : T648;
  assign T648 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_16;
  assign T649 = T557 & T650;
  assign T650 = T555[5'h10:5'h10];
  assign T967 = reset ? 1'h0 : T651;
  assign T651 = T653 ? 1'h1 : T652;
  assign T652 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_17;
  assign T653 = T557 & T654;
  assign T654 = T555[5'h11:5'h11];
  assign T655 = T556[1'h0:1'h0];
  assign T656 = T665 ? noCopyBaseAddr_19 : noCopyBaseAddr_18;
  assign T968 = reset ? 1'h0 : T657;
  assign T657 = T659 ? 1'h1 : T658;
  assign T658 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_18;
  assign T659 = T557 & T660;
  assign T660 = T555[5'h12:5'h12];
  assign T969 = reset ? 1'h0 : T661;
  assign T661 = T663 ? 1'h1 : T662;
  assign T662 = storeSeqMemConfig_io_rst ? 1'h0 : noCopyBaseAddr_19;
  assign T663 = T557 & T664;
  assign T664 = T555[5'h13:5'h13];
  assign T665 = T556[1'h0:1'h0];
  assign T666 = T556[1'h1:1'h1];
  assign T667 = T556[3'h4:3'h4];
  assign T668 = T970 + loopOffsetLkup;
  assign loopOffsetLkup = T669;
  assign T669 = T51 ? loopOffsetMem_io_outData : 32'h0;
  assign T970 = {23'h0, T672};
  assign T670 = T377 & T671;
  assign T671 = spillEndVal ^ 1'h1;
  assign T971 = {23'h0, T672};
  assign T792 = T544 & T793;
  assign T793 = T378 ^ 1'h1;
  assign T794 = baseAddrLkup - spillLkup;
  assign T795 = T796 & spillEndVal;
  assign T796 = T797 & T378;
  assign T797 = T51 & T798;
  assign T798 = noCopyBaseAddrVal ^ 1'h1;
  assign T799 = baseAddrLkup + loopOffsetLkup;
  assign T800 = T796 & T801;
  assign T801 = spillEndVal ^ 1'h1;
  assign baseAddrLkup = T802;
  assign T802 = T51 ? baseAddrMem_io_outData : 32'h0;
  assign T803 = T797 & T804;
  assign T804 = T378 ^ 1'h1;
  assign T805 = {storeReqAddr, storeReqData};
  assign T806 = {storeReqAddr, storeReqData};
  assign T807 = {storeReqAddr, storeReqData};
  assign T808 = {storeReqAddr, storeReqData};
  assign T809 = {storeReqAddr, storeReqData};
  assign T810 = {storeReqAddr, storeReqData};
  assign T811 = {storeReqAddr, storeReqData};
  assign T812 = {storeReqAddr, storeReqData};
  assign T813 = {storeReqAddr, storeReqData};
  assign T814 = {storeReqAddr, storeReqData};
  assign T815 = {storeReqAddr, storeReqData};
  assign T816 = {storeReqAddr, storeReqData};
  assign T817 = {storeReqAddr, storeReqData};
  assign T818 = {storeReqAddr, storeReqData};
  assign T819 = {storeReqAddr, storeReqData};
  assign T820 = {storeReqAddr, storeReqData};
  assign T821 = {storeReqAddr, storeReqData};
  assign T822 = {storeReqAddr, storeReqData};
  assign T823 = {storeReqAddr, storeReqData};
  assign T824 = T51 ? addrLkupIndex : 5'h0;
  assign T825 = T51 ? 1'h1 : 1'h0;
  assign T826 = T51 ? addrLkupIndex : 5'h0;
  assign T827 = T51 ? 1'h1 : 1'h0;
  assign T828 = io_seqMemAddrValid ? io_seqMemAddr : 9'h0;
  assign T829 = io_seqMemAddrValid ? io_seqMemAddrValid : 1'h0;
  assign T830 = T51 ? addrLkupIndex : 5'h0;
  assign T831 = T51 ? 1'h1 : 1'h0;
  assign io_computeDone = computeDone;
  assign computeDone = T832;
  assign T832 = T839 ? 1'h0 : T833;
  assign T833 = T834 & io_storeMemRdy;
  assign T834 = compDoneCnt == 3'h2;
  assign T972 = reset ? 3'h0 : T835;
  assign T835 = T838 ? T837 : T836;
  assign T836 = storeSeqMemConfig_io_rst ? 3'h0 : compDoneCnt;
  assign T837 = compDoneCnt + 3'h1;
  assign T838 = io_computeDoneCtrl & getNextReq;
  assign T839 = T833 ^ 1'h1;
  assign io_seqProceed = T840;
  assign T840 = T231 ? 1'h0 : T841;
  assign T841 = T225 ? 1'h1 : T842;
  assign T842 = T224 ? 1'h0 : T843;
  assign T843 = T218 ? 1'h1 : T844;
  assign T844 = T217 ? 1'h0 : T845;
  assign T845 = T211 ? 1'h1 : T846;
  assign T846 = T210 ? 1'h0 : T847;
  assign T847 = T204 ? 1'h1 : T848;
  assign T848 = T203 ? 1'h0 : T849;
  assign T849 = T197 ? 1'h1 : T850;
  assign T850 = T196 ? 1'h0 : T851;
  assign T851 = T190 ? 1'h1 : T852;
  assign T852 = T189 ? 1'h0 : T853;
  assign T853 = T183 ? 1'h1 : T854;
  assign T854 = T182 ? 1'h0 : T855;
  assign T855 = T176 ? 1'h1 : T856;
  assign T856 = T175 ? 1'h0 : T857;
  assign T857 = T169 ? 1'h1 : T858;
  assign T858 = T168 ? 1'h0 : T859;
  assign T859 = T162 ? 1'h1 : T860;
  assign T860 = T161 ? 1'h0 : T861;
  assign T861 = T155 ? 1'h1 : T862;
  assign T862 = T154 ? 1'h0 : T863;
  assign T863 = T148 ? 1'h1 : T864;
  assign T864 = T147 ? 1'h0 : T865;
  assign T865 = T141 ? 1'h1 : T866;
  assign T866 = T140 ? 1'h0 : T867;
  assign T867 = T134 ? 1'h1 : T868;
  assign T868 = T133 ? 1'h0 : T869;
  assign T869 = T127 ? 1'h1 : T870;
  assign T870 = T126 ? 1'h0 : T871;
  assign T871 = T120 ? 1'h1 : T872;
  assign T872 = T119 ? 1'h0 : T873;
  assign T873 = T113 ? 1'h1 : T874;
  assign T874 = T112 ? 1'h0 : T875;
  assign T875 = T106 ? 1'h1 : T876;
  assign T876 = T105 ? 1'h0 : T877;
  assign T877 = T99 ? 1'h1 : T878;
  assign T878 = T40 ? 1'h1 : 1'h0;
  assign io_storeMemValid = T879;
  assign T879 = io_storeMemRdy ? storeReqFifo_io_deqValid : 1'h0;
  assign io_storeMemData = T880;
  assign T880 = io_storeMemRdy ? storeReqFifo_io_deqData : 64'h0;
  customReg_1 baseAddrMem(.clk(clk),
       .io_inData( baseAddrMemConfig_io_memData ),
       .io_outData( baseAddrMem_io_outData ),
       .io_readEn( T831 ),
       .io_writeEn( baseAddrMemConfig_io_memOutValid ),
       .io_readAddr( T830 ),
       .io_writeAddr( baseAddrMemConfig_io_memAddr )
  );
  customReg_3 storeSeqMem(.clk(clk),
       .io_inData( storeSeqMemConfig_io_memData ),
       .io_outData( storeSeqMem_io_outData ),
       .io_readEn( T829 ),
       .io_writeEn( storeSeqMemConfig_io_memOutValid ),
       .io_readAddr( T828 ),
       .io_writeAddr( storeSeqMemConfig_io_memAddr )
  );
  customReg_1 loopOffsetMem(.clk(clk),
       .io_inData( loopOffsetMemConfig_io_memData ),
       .io_outData( loopOffsetMem_io_outData ),
       .io_readEn( T827 ),
       .io_writeEn( loopOffsetMemConfig_io_memOutValid ),
       .io_readAddr( T826 ),
       .io_writeAddr( loopOffsetMemConfig_io_memAddr )
  );
  customReg_1 spillOffsetMem(.clk(clk),
       .io_inData( spillOffsetMemConfig_io_memData ),
       .io_outData( spillOffsetMem_io_outData ),
       .io_readEn( T825 ),
       .io_writeEn( spillOffsetMemConfig_io_memOutValid ),
       .io_readAddr( T824 ),
       .io_writeAddr( spillOffsetMemConfig_io_memAddr )
  );
  memConfig_6 storeSeqMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( storeSeqMemConfig_io_memAddr ),
       .io_memData( storeSeqMemConfig_io_memData ),
       .io_memOutValid( storeSeqMemConfig_io_memOutValid ),
       .io_rst( storeSeqMemConfig_io_rst )
  );
  memConfig_7 baseAddrMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( baseAddrMemConfig_io_memAddr ),
       .io_memData( baseAddrMemConfig_io_memData ),
       .io_memOutValid( baseAddrMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  memConfig_8 loopOffsetMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( loopOffsetMemConfig_io_memAddr ),
       .io_memData( loopOffsetMemConfig_io_memData ),
       .io_memOutValid( loopOffsetMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  memConfig_9 spillOffsetMemConfig(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_memAddr( spillOffsetMemConfig_io_memAddr ),
       .io_memData( spillOffsetMemConfig_io_memData ),
       .io_memOutValid( spillOffsetMemConfig_io_memOutValid )
       //.io_rst(  )
  );
  fifo_5 storeReqFifo(.clk(clk), .reset(reset),
       .io_enqData( T233 ),
       .io_deqData( storeReqFifo_io_deqData ),
       .io_enqRdy( storeReqFifo_io_enqRdy ),
       .io_deqRdy( T232 ),
       .io_enqValid( T1 ),
       .io_deqValid( storeReqFifo_io_deqValid ),
       .io_rst( T0 )
  );

  always @(posedge clk) begin
    if(reset) begin
      portSel_0 <= 1'h0;
    end else if(T40) begin
      portSel_0 <= 1'h0;
    end else if(T44) begin
      portSel_0 <= 1'h1;
    end
    if(reset) begin
      nextSeq <= 43'h0;
    end else if(io_seqMemAddrValid) begin
      nextSeq <= storeSeqMem_io_outData;
    end
    if(reset) begin
      nextSeqValid <= 1'h0;
    end else if(T51) begin
      nextSeqValid <= 1'h0;
    end else if(storeSeqMemConfig_io_rst) begin
      nextSeqValid <= 1'h0;
    end else if(io_seqMemAddrValid) begin
      nextSeqValid <= 1'h1;
    end
    if(reset) begin
      firstReqDone <= 1'h0;
    end else if(T51) begin
      firstReqDone <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      firstReqDone <= 1'h0;
    end
    if(reset) begin
      portSel_1 <= 1'h0;
    end else if(T99) begin
      portSel_1 <= 1'h0;
    end else if(T103) begin
      portSel_1 <= 1'h1;
    end
    if(reset) begin
      portSel_2 <= 1'h0;
    end else if(T106) begin
      portSel_2 <= 1'h0;
    end else if(T110) begin
      portSel_2 <= 1'h1;
    end
    if(reset) begin
      portSel_3 <= 1'h0;
    end else if(T113) begin
      portSel_3 <= 1'h0;
    end else if(T117) begin
      portSel_3 <= 1'h1;
    end
    if(reset) begin
      portSel_4 <= 1'h0;
    end else if(T120) begin
      portSel_4 <= 1'h0;
    end else if(T124) begin
      portSel_4 <= 1'h1;
    end
    if(reset) begin
      portSel_5 <= 1'h0;
    end else if(T127) begin
      portSel_5 <= 1'h0;
    end else if(T131) begin
      portSel_5 <= 1'h1;
    end
    if(reset) begin
      portSel_6 <= 1'h0;
    end else if(T134) begin
      portSel_6 <= 1'h0;
    end else if(T138) begin
      portSel_6 <= 1'h1;
    end
    if(reset) begin
      portSel_7 <= 1'h0;
    end else if(T141) begin
      portSel_7 <= 1'h0;
    end else if(T145) begin
      portSel_7 <= 1'h1;
    end
    if(reset) begin
      portSel_8 <= 1'h0;
    end else if(T148) begin
      portSel_8 <= 1'h0;
    end else if(T152) begin
      portSel_8 <= 1'h1;
    end
    if(reset) begin
      portSel_9 <= 1'h0;
    end else if(T155) begin
      portSel_9 <= 1'h0;
    end else if(T159) begin
      portSel_9 <= 1'h1;
    end
    if(reset) begin
      portSel_10 <= 1'h0;
    end else if(T162) begin
      portSel_10 <= 1'h0;
    end else if(T166) begin
      portSel_10 <= 1'h1;
    end
    if(reset) begin
      portSel_11 <= 1'h0;
    end else if(T169) begin
      portSel_11 <= 1'h0;
    end else if(T173) begin
      portSel_11 <= 1'h1;
    end
    if(reset) begin
      portSel_12 <= 1'h0;
    end else if(T176) begin
      portSel_12 <= 1'h0;
    end else if(T180) begin
      portSel_12 <= 1'h1;
    end
    if(reset) begin
      portSel_13 <= 1'h0;
    end else if(T183) begin
      portSel_13 <= 1'h0;
    end else if(T187) begin
      portSel_13 <= 1'h1;
    end
    if(reset) begin
      portSel_14 <= 1'h0;
    end else if(T190) begin
      portSel_14 <= 1'h0;
    end else if(T194) begin
      portSel_14 <= 1'h1;
    end
    if(reset) begin
      portSel_15 <= 1'h0;
    end else if(T197) begin
      portSel_15 <= 1'h0;
    end else if(T201) begin
      portSel_15 <= 1'h1;
    end
    if(reset) begin
      portSel_16 <= 1'h0;
    end else if(T204) begin
      portSel_16 <= 1'h0;
    end else if(T208) begin
      portSel_16 <= 1'h1;
    end
    if(reset) begin
      portSel_17 <= 1'h0;
    end else if(T211) begin
      portSel_17 <= 1'h0;
    end else if(T215) begin
      portSel_17 <= 1'h1;
    end
    if(reset) begin
      portSel_18 <= 1'h0;
    end else if(T218) begin
      portSel_18 <= 1'h0;
    end else if(T222) begin
      portSel_18 <= 1'h1;
    end
    if(reset) begin
      portSel_19 <= 1'h0;
    end else if(T225) begin
      portSel_19 <= 1'h0;
    end else if(T229) begin
      portSel_19 <= 1'h1;
    end
    if(reset) begin
      storeMemAddr <= 32'h0;
    end else if(T51) begin
      storeMemAddr <= T354;
    end
    if(reset) begin
      savedOffsets_0 <= 9'h0;
    end else if(T679) begin
      savedOffsets_0 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_0 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_1 <= 9'h0;
    end else if(T685) begin
      savedOffsets_1 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_1 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_2 <= 9'h0;
    end else if(T691) begin
      savedOffsets_2 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_2 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_3 <= 9'h0;
    end else if(T695) begin
      savedOffsets_3 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_3 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_4 <= 9'h0;
    end else if(T703) begin
      savedOffsets_4 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_4 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_5 <= 9'h0;
    end else if(T707) begin
      savedOffsets_5 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_5 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_6 <= 9'h0;
    end else if(T713) begin
      savedOffsets_6 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_6 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_7 <= 9'h0;
    end else if(T717) begin
      savedOffsets_7 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_7 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_8 <= 9'h0;
    end else if(T727) begin
      savedOffsets_8 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_8 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_9 <= 9'h0;
    end else if(T731) begin
      savedOffsets_9 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_9 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_10 <= 9'h0;
    end else if(T737) begin
      savedOffsets_10 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_10 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_11 <= 9'h0;
    end else if(T741) begin
      savedOffsets_11 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_11 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_12 <= 9'h0;
    end else if(T749) begin
      savedOffsets_12 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_12 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_13 <= 9'h0;
    end else if(T753) begin
      savedOffsets_13 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_13 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_14 <= 9'h0;
    end else if(T759) begin
      savedOffsets_14 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_14 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_15 <= 9'h0;
    end else if(T763) begin
      savedOffsets_15 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_15 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_16 <= 9'h0;
    end else if(T773) begin
      savedOffsets_16 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_16 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_17 <= 9'h0;
    end else if(T777) begin
      savedOffsets_17 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_17 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_18 <= 9'h0;
    end else if(T783) begin
      savedOffsets_18 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_18 <= 9'h0;
    end
    if(reset) begin
      savedOffsets_19 <= 9'h0;
    end else if(T787) begin
      savedOffsets_19 <= savedOffsetsVal;
    end else if(storeSeqMemConfig_io_rst) begin
      savedOffsets_19 <= 9'h0;
    end
    if(reset) begin
      spillEnd <= 1'h0;
    end else if(storeSeqMemConfig_io_rst) begin
      spillEnd <= 1'h0;
    end else if(io_seqMemAddrValid) begin
      spillEnd <= io_spillEnd;
    end
    if(reset) begin
      nextIterStart <= 1'h0;
    end else if(io_seqMemAddrValid) begin
      nextIterStart <= io_nextIterStart;
    end
    if(reset) begin
      offsetUpdate_0 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_0 <= offsetUpdateVal_0;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_0 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_1 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_1 <= offsetUpdateVal_1;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_1 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_2 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_2 <= offsetUpdateVal_2;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_2 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_3 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_3 <= offsetUpdateVal_3;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_3 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_4 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_4 <= offsetUpdateVal_4;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_4 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_5 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_5 <= offsetUpdateVal_5;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_5 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_6 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_6 <= offsetUpdateVal_6;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_6 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_7 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_7 <= offsetUpdateVal_7;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_7 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_8 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_8 <= offsetUpdateVal_8;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_8 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_9 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_9 <= offsetUpdateVal_9;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_9 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_10 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_10 <= offsetUpdateVal_10;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_10 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_11 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_11 <= offsetUpdateVal_11;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_11 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_12 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_12 <= offsetUpdateVal_12;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_12 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_13 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_13 <= offsetUpdateVal_13;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_13 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_14 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_14 <= offsetUpdateVal_14;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_14 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_15 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_15 <= offsetUpdateVal_15;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_15 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_16 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_16 <= offsetUpdateVal_16;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_16 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_17 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_17 <= offsetUpdateVal_17;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_17 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_18 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_18 <= offsetUpdateVal_18;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_18 <= 1'h0;
    end
    if(reset) begin
      offsetUpdate_19 <= 1'h0;
    end else if(T51) begin
      offsetUpdate_19 <= offsetUpdateVal_19;
    end else if(storeSeqMemConfig_io_rst) begin
      offsetUpdate_19 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_0 <= 1'h0;
    end else if(T553) begin
      noCopyBaseAddr_0 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_0 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_1 <= 1'h0;
    end else if(T561) begin
      noCopyBaseAddr_1 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_1 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_2 <= 1'h0;
    end else if(T567) begin
      noCopyBaseAddr_2 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_2 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_3 <= 1'h0;
    end else if(T571) begin
      noCopyBaseAddr_3 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_3 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_4 <= 1'h0;
    end else if(T579) begin
      noCopyBaseAddr_4 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_4 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_5 <= 1'h0;
    end else if(T583) begin
      noCopyBaseAddr_5 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_5 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_6 <= 1'h0;
    end else if(T589) begin
      noCopyBaseAddr_6 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_6 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_7 <= 1'h0;
    end else if(T593) begin
      noCopyBaseAddr_7 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_7 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_8 <= 1'h0;
    end else if(T603) begin
      noCopyBaseAddr_8 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_8 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_9 <= 1'h0;
    end else if(T607) begin
      noCopyBaseAddr_9 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_9 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_10 <= 1'h0;
    end else if(T613) begin
      noCopyBaseAddr_10 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_10 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_11 <= 1'h0;
    end else if(T617) begin
      noCopyBaseAddr_11 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_11 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_12 <= 1'h0;
    end else if(T625) begin
      noCopyBaseAddr_12 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_12 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_13 <= 1'h0;
    end else if(T629) begin
      noCopyBaseAddr_13 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_13 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_14 <= 1'h0;
    end else if(T635) begin
      noCopyBaseAddr_14 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_14 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_15 <= 1'h0;
    end else if(T639) begin
      noCopyBaseAddr_15 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_15 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_16 <= 1'h0;
    end else if(T649) begin
      noCopyBaseAddr_16 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_16 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_17 <= 1'h0;
    end else if(T653) begin
      noCopyBaseAddr_17 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_17 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_18 <= 1'h0;
    end else if(T659) begin
      noCopyBaseAddr_18 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_18 <= 1'h0;
    end
    if(reset) begin
      noCopyBaseAddr_19 <= 1'h0;
    end else if(T663) begin
      noCopyBaseAddr_19 <= 1'h1;
    end else if(storeSeqMemConfig_io_rst) begin
      noCopyBaseAddr_19 <= 1'h0;
    end
    if(reset) begin
      compDoneCnt <= 3'h0;
    end else if(T838) begin
      compDoneCnt <= T837;
    end else if(storeSeqMemConfig_io_rst) begin
      compDoneCnt <= 3'h0;
    end
  end
endmodule

module storeSeq(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    input [31:0] io_fabOutToStore_19,
    input [31:0] io_fabOutToStore_18,
    input [31:0] io_fabOutToStore_17,
    input [31:0] io_fabOutToStore_16,
    input [31:0] io_fabOutToStore_15,
    input [31:0] io_fabOutToStore_14,
    input [31:0] io_fabOutToStore_13,
    input [31:0] io_fabOutToStore_12,
    input [31:0] io_fabOutToStore_11,
    input [31:0] io_fabOutToStore_10,
    input [31:0] io_fabOutToStore_9,
    input [31:0] io_fabOutToStore_8,
    input [31:0] io_fabOutToStore_7,
    input [31:0] io_fabOutToStore_6,
    input [31:0] io_fabOutToStore_5,
    input [31:0] io_fabOutToStore_4,
    input [31:0] io_fabOutToStore_3,
    input [31:0] io_fabOutToStore_2,
    input [31:0] io_fabOutToStore_1,
    input [31:0] io_fabOutToStore_0,
    input  io_fabOutToStoreValid_19,
    input  io_fabOutToStoreValid_18,
    input  io_fabOutToStoreValid_17,
    input  io_fabOutToStoreValid_16,
    input  io_fabOutToStoreValid_15,
    input  io_fabOutToStoreValid_14,
    input  io_fabOutToStoreValid_13,
    input  io_fabOutToStoreValid_12,
    input  io_fabOutToStoreValid_11,
    input  io_fabOutToStoreValid_10,
    input  io_fabOutToStoreValid_9,
    input  io_fabOutToStoreValid_8,
    input  io_fabOutToStoreValid_7,
    input  io_fabOutToStoreValid_6,
    input  io_fabOutToStoreValid_5,
    input  io_fabOutToStoreValid_4,
    input  io_fabOutToStoreValid_3,
    input  io_fabOutToStoreValid_2,
    input  io_fabOutToStoreValid_1,
    input  io_fabOutToStoreValid_0,
    output[63:0] io_storeMemData,
    output io_storeMemValid,
    input  io_storeMemRdy,
    output io_computeDone
);

  wire storeCtrlClass_io_spillEnd;
  wire storeCtrlClass_io_nextIterStart;
  wire[8:0] storeCtrlClass_io_seqMemAddr;
  wire storeCtrlClass_io_seqMemAddrValid;
  wire storeCtrlClass_io_computeDone;
  wire[63:0] storeDPClass_io_storeMemData;
  wire storeDPClass_io_storeMemValid;
  wire storeDPClass_io_seqProceed;
  wire storeDPClass_io_computeDone;


  assign io_computeDone = storeDPClass_io_computeDone;
  assign io_storeMemValid = storeDPClass_io_storeMemValid;
  assign io_storeMemData = storeDPClass_io_storeMemData;
  storeSeqCtrl storeCtrlClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_spillEnd( storeCtrlClass_io_spillEnd ),
       .io_nextIterStart( storeCtrlClass_io_nextIterStart ),
       .io_seqMemAddr( storeCtrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( storeCtrlClass_io_seqMemAddrValid ),
       .io_seqProceed( storeDPClass_io_seqProceed ),
       .io_computeDone( storeCtrlClass_io_computeDone )
  );
  storeSeqDP storeDPClass(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       .io_inValid( io_inValid ),
       .io_spillEnd( storeCtrlClass_io_spillEnd ),
       .io_nextIterStart( storeCtrlClass_io_nextIterStart ),
       .io_seqMemAddr( storeCtrlClass_io_seqMemAddr ),
       .io_seqMemAddrValid( storeCtrlClass_io_seqMemAddrValid ),
       .io_storeMemData( storeDPClass_io_storeMemData ),
       .io_storeMemValid( storeDPClass_io_storeMemValid ),
       .io_storeMemRdy( io_storeMemRdy ),
       .io_seqProceed( storeDPClass_io_seqProceed ),
       .io_fabOutToStore_19( io_fabOutToStore_19 ),
       .io_fabOutToStore_18( io_fabOutToStore_18 ),
       .io_fabOutToStore_17( io_fabOutToStore_17 ),
       .io_fabOutToStore_16( io_fabOutToStore_16 ),
       .io_fabOutToStore_15( io_fabOutToStore_15 ),
       .io_fabOutToStore_14( io_fabOutToStore_14 ),
       .io_fabOutToStore_13( io_fabOutToStore_13 ),
       .io_fabOutToStore_12( io_fabOutToStore_12 ),
       .io_fabOutToStore_11( io_fabOutToStore_11 ),
       .io_fabOutToStore_10( io_fabOutToStore_10 ),
       .io_fabOutToStore_9( io_fabOutToStore_9 ),
       .io_fabOutToStore_8( io_fabOutToStore_8 ),
       .io_fabOutToStore_7( io_fabOutToStore_7 ),
       .io_fabOutToStore_6( io_fabOutToStore_6 ),
       .io_fabOutToStore_5( io_fabOutToStore_5 ),
       .io_fabOutToStore_4( io_fabOutToStore_4 ),
       .io_fabOutToStore_3( io_fabOutToStore_3 ),
       .io_fabOutToStore_2( io_fabOutToStore_2 ),
       .io_fabOutToStore_1( io_fabOutToStore_1 ),
       .io_fabOutToStore_0( io_fabOutToStore_0 ),
       .io_fabOutToStoreValid_19( io_fabOutToStoreValid_19 ),
       .io_fabOutToStoreValid_18( io_fabOutToStoreValid_18 ),
       .io_fabOutToStoreValid_17( io_fabOutToStoreValid_17 ),
       .io_fabOutToStoreValid_16( io_fabOutToStoreValid_16 ),
       .io_fabOutToStoreValid_15( io_fabOutToStoreValid_15 ),
       .io_fabOutToStoreValid_14( io_fabOutToStoreValid_14 ),
       .io_fabOutToStoreValid_13( io_fabOutToStoreValid_13 ),
       .io_fabOutToStoreValid_12( io_fabOutToStoreValid_12 ),
       .io_fabOutToStoreValid_11( io_fabOutToStoreValid_11 ),
       .io_fabOutToStoreValid_10( io_fabOutToStoreValid_10 ),
       .io_fabOutToStoreValid_9( io_fabOutToStoreValid_9 ),
       .io_fabOutToStoreValid_8( io_fabOutToStoreValid_8 ),
       .io_fabOutToStoreValid_7( io_fabOutToStoreValid_7 ),
       .io_fabOutToStoreValid_6( io_fabOutToStoreValid_6 ),
       .io_fabOutToStoreValid_5( io_fabOutToStoreValid_5 ),
       .io_fabOutToStoreValid_4( io_fabOutToStoreValid_4 ),
       .io_fabOutToStoreValid_3( io_fabOutToStoreValid_3 ),
       .io_fabOutToStoreValid_2( io_fabOutToStoreValid_2 ),
       .io_fabOutToStoreValid_1( io_fabOutToStoreValid_1 ),
       .io_fabOutToStoreValid_0( io_fabOutToStoreValid_0 ),
       .io_computeDone( storeDPClass_io_computeDone ),
       .io_computeDoneCtrl( storeCtrlClass_io_computeDone )
  );
endmodule

module mainConfigure(input clk, input reset,
    input [31:0] io_configData,
    input  io_configDataValid,
    output[31:0] io_loadConfig,
    output io_loadConfigValid,
    output[31:0] io_storeConfig,
    output io_storeConfigValid,
    output[31:0] io_fabInConfig,
    output io_fabInConfigValid,
    output[31:0] io_fabOutConfig,
    output io_fabOutConfigValid,
    output[31:0] io_fabConfig,
    output io_fabConfigValid
);

  reg  configValidReg;
  wire T0;
  reg [31:0] configReg;
  wire[31:0] T1;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    configValidReg = {1{$random}};
    configReg = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign io_loadConfigValid = {1{$random}};
  assign io_loadConfig = {1{$random}};
// synthesis translate_on
`endif
  assign io_fabConfigValid = configValidReg;
  assign T0 = reset ? 1'h0 : io_configDataValid;
  assign io_fabConfig = configReg;
  assign T1 = reset ? 32'h0 : io_configData;
  assign io_fabOutConfigValid = configValidReg;
  assign io_fabOutConfig = configReg;
  assign io_fabInConfigValid = configValidReg;
  assign io_fabInConfig = configReg;
  assign io_storeConfigValid = configValidReg;
  assign io_storeConfig = configReg;

  always @(posedge clk) begin
    if(reset) begin
      configValidReg <= 1'h0;
    end else begin
      configValidReg <= io_configDataValid;
    end
    if(reset) begin
      configReg <= 32'h0;
    end else begin
      configReg <= io_configData;
    end
  end
endmodule

module fabricConfigure_0(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h0;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigure_1(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h1;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigure_2(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h2;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigure_3(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h3;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigure_4(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h4;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigure_5(input clk, input reset,
    input [31:0] io_inConfig,
    //input  io_inValid
    output[32:0] io_outConfig,
    //output io_outValid
    input  io_rst
);

  reg [32:0] outDataReg;
  wire[32:0] T93;
  wire[32:0] T0;
  wire[32:0] T1;
  wire[32:0] T2;
  wire[32:0] T3;
  wire[32:0] T4;
  wire[32:0] T5;
  wire[32:0] T6;
  wire[32:0] T7;
  wire[32:0] T8;
  wire[32:0] T9;
  wire[32:0] T10;
  wire[32:0] T11;
  wire[32:0] T94;
  wire T12;
  wire T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[32:0] T16;
  wire[32:0] T95;
  wire[31:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [31:0] inDataReg;
  wire[31:0] T96;
  wire[32:0] T20;
  wire[32:0] T21;
  wire[32:0] T22;
  wire[32:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  configValid;
  wire T97;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[2:0] ownIndex;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[32:0] T46;
  wire[32:0] T47;
  wire[32:0] T48;
  wire[32:0] T49;
  wire[32:0] T98;
  wire T50;
  wire T51;
  wire[32:0] T52;
  wire[32:0] T53;
  wire[32:0] T54;
  wire[32:0] T55;
  wire[32:0] T56;
  wire[32:0] T57;
  wire[32:0] T58;
  wire[32:0] T59;
  wire[32:0] T99;
  wire[12:0] T60;
  wire[12:0] T61;
  wire[12:0] T62;
  wire[32:0] T63;
  wire[32:0] T64;
  wire[32:0] T65;
  wire[32:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[32:0] T70;
  wire[32:0] T71;
  wire[32:0] T72;
  wire[32:0] T73;
  wire[32:0] T100;
  wire T74;
  wire T75;
  wire[32:0] T76;
  wire[32:0] T77;
  wire[32:0] T78;
  wire[32:0] T79;
  wire[32:0] T80;
  wire[32:0] T81;
  wire[32:0] T82;
  wire[32:0] T83;
  wire[32:0] T101;
  wire[23:0] T84;
  wire[23:0] T85;
  wire[23:0] T86;
  wire[32:0] T87;
  wire[32:0] T88;
  wire[32:0] T89;
  wire[32:0] T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    outDataReg = {2{$random}};
    inDataReg = {1{$random}};
    configValid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_outValid = {1{$random}};
// synthesis translate_on
`endif
  assign io_outConfig = outDataReg;
  assign T93 = reset ? 33'h0 : T0;
  assign T0 = T91 ? T83 : T1;
  assign T1 = T91 ? T78 : T2;
  assign T2 = T91 ? T70 : T3;
  assign T3 = T67 ? T59 : T4;
  assign T4 = T67 ? T54 : T5;
  assign T5 = T67 ? T46 : T6;
  assign T6 = T24 ? T16 : T7;
  assign T7 = T24 ? T8 : outDataReg;
  assign T8 = T14 | T9;
  assign T9 = T94 & T10;
  assign T10 = 33'h100000000 | T11;
  assign T11 = outDataReg ^ outDataReg;
  assign T94 = T12 ? 33'h1ffffffff : 33'h0;
  assign T12 = T13;
  assign T13 = 1'h1;
  assign T14 = outDataReg & T15;
  assign T15 = ~ T10;
  assign T16 = T20 | T95;
  assign T95 = {1'h0, T17};
  assign T17 = T18 << 5'h1d;
  assign T18 = T19 & 3'h7;
  assign T19 = inDataReg[5'h1b:5'h19];
  assign T96 = reset ? 32'h0 : io_inConfig;
  assign T20 = T7 & T21;
  assign T21 = ~ T22;
  assign T22 = 33'he0000000 | T23;
  assign T23 = outDataReg ^ outDataReg;
  assign T24 = T27 & T25;
  assign T25 = T26 == 2'h1;
  assign T26 = inDataReg[5'h1e:5'h1d];
  assign T27 = T44 & configValid;
  assign T97 = reset ? 1'h0 : T28;
  assign T28 = io_rst ? 1'h0 : T29;
  assign T29 = T42 ? 1'h0 : T30;
  assign T30 = T40 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : configValid;
  assign T32 = T35 & T33;
  assign T33 = T34 == ownIndex;
  assign ownIndex = 3'h5;
  assign T34 = inDataReg[2'h2:1'h0];
  assign T35 = T38 & T36;
  assign T36 = T37 == 2'h1;
  assign T37 = inDataReg[5'h1e:5'h1d];
  assign T38 = T39 == 1'h0;
  assign T39 = inDataReg[5'h1f:5'h1f];
  assign T40 = T35 & T41;
  assign T41 = T33 ^ 1'h1;
  assign T42 = T38 & T43;
  assign T43 = T36 ^ 1'h1;
  assign T44 = T45 == 1'h1;
  assign T45 = inDataReg[5'h1f:5'h1f];
  assign T46 = T52 | T47;
  assign T47 = T98 & T48;
  assign T48 = 33'h10000000 | T49;
  assign T49 = outDataReg ^ outDataReg;
  assign T98 = T50 ? 33'h1ffffffff : 33'h0;
  assign T50 = T51;
  assign T51 = 1'h0;
  assign T52 = T6 & T53;
  assign T53 = ~ T48;
  assign T54 = T55 | 33'h0;
  assign T55 = T5 & T56;
  assign T56 = ~ T57;
  assign T57 = 33'hfffe000 | T58;
  assign T58 = outDataReg ^ outDataReg;
  assign T59 = T63 | T99;
  assign T99 = {20'h0, T60};
  assign T60 = T61 << 1'h0;
  assign T61 = T62 & 13'h1fff;
  assign T62 = inDataReg[4'hc:1'h0];
  assign T63 = T4 & T64;
  assign T64 = ~ T65;
  assign T65 = 33'h1fff | T66;
  assign T66 = outDataReg ^ outDataReg;
  assign T67 = T24 & T68;
  assign T68 = T69;
  assign T69 = inDataReg[5'h18:5'h18];
  assign T70 = T76 | T71;
  assign T71 = T100 & T72;
  assign T72 = 33'h10000000 | T73;
  assign T73 = outDataReg ^ outDataReg;
  assign T100 = T74 ? 33'h1ffffffff : 33'h0;
  assign T74 = T75;
  assign T75 = 1'h1;
  assign T76 = T3 & T77;
  assign T77 = ~ T72;
  assign T78 = T79 | 33'h0;
  assign T79 = T2 & T80;
  assign T80 = ~ T81;
  assign T81 = 33'hf000000 | T82;
  assign T82 = outDataReg ^ outDataReg;
  assign T83 = T87 | T101;
  assign T101 = {9'h0, T84};
  assign T84 = T85 << 1'h0;
  assign T85 = T86 & 24'hffffff;
  assign T86 = inDataReg[5'h17:1'h0];
  assign T87 = T1 & T88;
  assign T88 = ~ T89;
  assign T89 = 33'hffffff | T90;
  assign T90 = outDataReg ^ outDataReg;
  assign T91 = T24 & T92;
  assign T92 = T68 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      outDataReg <= 33'h0;
    end else if(T91) begin
      outDataReg <= T83;
    end else if(T91) begin
      outDataReg <= T78;
    end else if(T91) begin
      outDataReg <= T70;
    end else if(T67) begin
      outDataReg <= T59;
    end else if(T67) begin
      outDataReg <= T54;
    end else if(T67) begin
      outDataReg <= T46;
    end else if(T24) begin
      outDataReg <= T16;
    end else if(T24) begin
      outDataReg <= T8;
    end
    if(reset) begin
      inDataReg <= 32'h0;
    end else begin
      inDataReg <= io_inConfig;
    end
    if(reset) begin
      configValid <= 1'h0;
    end else if(io_rst) begin
      configValid <= 1'h0;
    end else if(T42) begin
      configValid <= 1'h0;
    end else if(T40) begin
      configValid <= 1'h0;
    end else if(T32) begin
      configValid <= 1'h1;
    end
  end
endmodule

module fabricConfigureTop(input clk, input reset,
    input [31:0] io_inConfig,
    output[32:0] io_outConfig_5,
    output[32:0] io_outConfig_4,
    output[32:0] io_outConfig_3,
    output[32:0] io_outConfig_2,
    output[32:0] io_outConfig_1,
    output[32:0] io_outConfig_0,
    input  io_rst
);

  wire[32:0] fabricConfigure_io_outConfig;
  wire[32:0] fabricConfigure_1_io_outConfig;
  wire[32:0] fabricConfigure_2_io_outConfig;
  wire[32:0] fabricConfigure_3_io_outConfig;
  wire[32:0] fabricConfigure_4_io_outConfig;
  wire[32:0] fabricConfigure_5_io_outConfig;


  assign io_outConfig_0 = fabricConfigure_io_outConfig;
  assign io_outConfig_1 = fabricConfigure_1_io_outConfig;
  assign io_outConfig_2 = fabricConfigure_2_io_outConfig;
  assign io_outConfig_3 = fabricConfigure_3_io_outConfig;
  assign io_outConfig_4 = fabricConfigure_4_io_outConfig;
  assign io_outConfig_5 = fabricConfigure_5_io_outConfig;
  fabricConfigure_0 fabricConfigure(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
  fabricConfigure_1 fabricConfigure_1(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_1_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
  fabricConfigure_2 fabricConfigure_2(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_2_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
  fabricConfigure_3 fabricConfigure_3(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_3_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
  fabricConfigure_4 fabricConfigure_4(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_4_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
  fabricConfigure_5 fabricConfigure_5(.clk(clk), .reset(reset),
       .io_inConfig( io_inConfig ),
       //.io_inValid(  )
       .io_outConfig( fabricConfigure_5_io_outConfig ),
       //.io_outValid(  )
       .io_rst( io_rst )
  );
endmodule

module controllerTop(input clk, input reset,
    input [31:0] io_inConfig,
    input  io_inValid,
    output[31:0] io_loadRqst,
    output io_loadRqstValid,
    input  io_loadRqstRdy,
    input [37:0] io_loadResp,
    input  io_loadRespValid,
    output io_loadRespRdy,
    output[63:0] io_storeMemData,
    output io_storeMemValid,
    input  io_storeMemRdy,
    output[31:0] io_fabInData_19,
    output[31:0] io_fabInData_18,
    output[31:0] io_fabInData_17,
    output[31:0] io_fabInData_16,
    output[31:0] io_fabInData_15,
    output[31:0] io_fabInData_14,
    output[31:0] io_fabInData_13,
    output[31:0] io_fabInData_12,
    output[31:0] io_fabInData_11,
    output[31:0] io_fabInData_10,
    output[31:0] io_fabInData_9,
    output[31:0] io_fabInData_8,
    output[31:0] io_fabInData_7,
    output[31:0] io_fabInData_6,
    output[31:0] io_fabInData_5,
    output[31:0] io_fabInData_4,
    output[31:0] io_fabInData_3,
    output[31:0] io_fabInData_2,
    output[31:0] io_fabInData_1,
    output[31:0] io_fabInData_0,
    output io_fabInValid_19,
    output io_fabInValid_18,
    output io_fabInValid_17,
    output io_fabInValid_16,
    output io_fabInValid_15,
    output io_fabInValid_14,
    output io_fabInValid_13,
    output io_fabInValid_12,
    output io_fabInValid_11,
    output io_fabInValid_10,
    output io_fabInValid_9,
    output io_fabInValid_8,
    output io_fabInValid_7,
    output io_fabInValid_6,
    output io_fabInValid_5,
    output io_fabInValid_4,
    output io_fabInValid_3,
    output io_fabInValid_2,
    output io_fabInValid_1,
    output io_fabInValid_0,
    input  io_fabInRdy_19,
    input  io_fabInRdy_18,
    input  io_fabInRdy_17,
    input  io_fabInRdy_16,
    input  io_fabInRdy_15,
    input  io_fabInRdy_14,
    input  io_fabInRdy_13,
    input  io_fabInRdy_12,
    input  io_fabInRdy_11,
    input  io_fabInRdy_10,
    input  io_fabInRdy_9,
    input  io_fabInRdy_8,
    input  io_fabInRdy_7,
    input  io_fabInRdy_6,
    input  io_fabInRdy_5,
    input  io_fabInRdy_4,
    input  io_fabInRdy_3,
    input  io_fabInRdy_2,
    input  io_fabInRdy_1,
    input  io_fabInRdy_0,
    input [31:0] io_fabOut_19,
    input [31:0] io_fabOut_18,
    input [31:0] io_fabOut_17,
    input [31:0] io_fabOut_16,
    input [31:0] io_fabOut_15,
    input [31:0] io_fabOut_14,
    input [31:0] io_fabOut_13,
    input [31:0] io_fabOut_12,
    input [31:0] io_fabOut_11,
    input [31:0] io_fabOut_10,
    input [31:0] io_fabOut_9,
    input [31:0] io_fabOut_8,
    input [31:0] io_fabOut_7,
    input [31:0] io_fabOut_6,
    input [31:0] io_fabOut_5,
    input [31:0] io_fabOut_4,
    input [31:0] io_fabOut_3,
    input [31:0] io_fabOut_2,
    input [31:0] io_fabOut_1,
    input [31:0] io_fabOut_0,
    input  io_fabOutValid_19,
    input  io_fabOutValid_18,
    input  io_fabOutValid_17,
    input  io_fabOutValid_16,
    input  io_fabOutValid_15,
    input  io_fabOutValid_14,
    input  io_fabOutValid_13,
    input  io_fabOutValid_12,
    input  io_fabOutValid_11,
    input  io_fabOutValid_10,
    input  io_fabOutValid_9,
    input  io_fabOutValid_8,
    input  io_fabOutValid_7,
    input  io_fabOutValid_6,
    input  io_fabOutValid_5,
    input  io_fabOutValid_4,
    input  io_fabOutValid_3,
    input  io_fabOutValid_2,
    input  io_fabOutValid_1,
    input  io_fabOutValid_0,
    output io_fabOutRdy_19,
    output io_fabOutRdy_18,
    output io_fabOutRdy_17,
    output io_fabOutRdy_16,
    output io_fabOutRdy_15,
    output io_fabOutRdy_14,
    output io_fabOutRdy_13,
    output io_fabOutRdy_12,
    output io_fabOutRdy_11,
    output io_fabOutRdy_10,
    output io_fabOutRdy_9,
    output io_fabOutRdy_8,
    output io_fabOutRdy_7,
    output io_fabOutRdy_6,
    output io_fabOutRdy_5,
    output io_fabOutRdy_4,
    output io_fabOutRdy_3,
    output io_fabOutRdy_2,
    output io_fabOutRdy_1,
    output io_fabOutRdy_0
);

  wire[37:0] T0;
  wire[37:0] T1;
  wire[37:0] T2;
  wire[37:0] T3;
  wire[37:0] T4;
  wire[37:0] T5;
  wire[37:0] T6;
  wire[37:0] T7;
  wire[31:0] mainConfigClass_io_loadConfig;
  wire mainConfigClass_io_loadConfigValid;
  wire[31:0] mainConfigClass_io_storeConfig;
  wire mainConfigClass_io_storeConfigValid;
  wire[31:0] mainConfigClass_io_fabInConfig;
  wire mainConfigClass_io_fabInConfigValid;
  wire[31:0] mainConfigClass_io_fabOutConfig;
  wire mainConfigClass_io_fabOutConfigValid;
  wire[31:0] loadSeqClass_io_loadRqst;
  wire loadSeqClass_io_loadRqstValid;
  wire loadSeqClass_io_loadRespRdy;
  wire[37:0] loadSeqClass_io_memBankEnq_7;
  wire[37:0] loadSeqClass_io_memBankEnq_6;
  wire[37:0] loadSeqClass_io_memBankEnq_5;
  wire[37:0] loadSeqClass_io_memBankEnq_4;
  wire[37:0] loadSeqClass_io_memBankEnq_3;
  wire[37:0] loadSeqClass_io_memBankEnq_2;
  wire[37:0] loadSeqClass_io_memBankEnq_1;
  wire[37:0] loadSeqClass_io_memBankEnq_0;
  wire loadSeqClass_io_memBankValid_7;
  wire loadSeqClass_io_memBankValid_6;
  wire loadSeqClass_io_memBankValid_5;
  wire loadSeqClass_io_memBankValid_4;
  wire loadSeqClass_io_memBankValid_3;
  wire loadSeqClass_io_memBankValid_2;
  wire loadSeqClass_io_memBankValid_1;
  wire loadSeqClass_io_memBankValid_0;
  wire[63:0] storeSeqClass_io_storeMemData;
  wire storeSeqClass_io_storeMemValid;
  wire fabOutSeqClass_io_fabOutRdy_19;
  wire fabOutSeqClass_io_fabOutRdy_18;
  wire fabOutSeqClass_io_fabOutRdy_17;
  wire fabOutSeqClass_io_fabOutRdy_16;
  wire fabOutSeqClass_io_fabOutRdy_15;
  wire fabOutSeqClass_io_fabOutRdy_14;
  wire fabOutSeqClass_io_fabOutRdy_13;
  wire fabOutSeqClass_io_fabOutRdy_12;
  wire fabOutSeqClass_io_fabOutRdy_11;
  wire fabOutSeqClass_io_fabOutRdy_10;
  wire fabOutSeqClass_io_fabOutRdy_9;
  wire fabOutSeqClass_io_fabOutRdy_8;
  wire fabOutSeqClass_io_fabOutRdy_7;
  wire fabOutSeqClass_io_fabOutRdy_6;
  wire fabOutSeqClass_io_fabOutRdy_5;
  wire fabOutSeqClass_io_fabOutRdy_4;
  wire fabOutSeqClass_io_fabOutRdy_3;
  wire fabOutSeqClass_io_fabOutRdy_2;
  wire fabOutSeqClass_io_fabOutRdy_1;
  wire fabOutSeqClass_io_fabOutRdy_0;
  wire[31:0] fabOutSeqClass_io_fabOutStore_19;
  wire[31:0] fabOutSeqClass_io_fabOutStore_18;
  wire[31:0] fabOutSeqClass_io_fabOutStore_17;
  wire[31:0] fabOutSeqClass_io_fabOutStore_16;
  wire[31:0] fabOutSeqClass_io_fabOutStore_15;
  wire[31:0] fabOutSeqClass_io_fabOutStore_14;
  wire[31:0] fabOutSeqClass_io_fabOutStore_13;
  wire[31:0] fabOutSeqClass_io_fabOutStore_12;
  wire[31:0] fabOutSeqClass_io_fabOutStore_11;
  wire[31:0] fabOutSeqClass_io_fabOutStore_10;
  wire[31:0] fabOutSeqClass_io_fabOutStore_9;
  wire[31:0] fabOutSeqClass_io_fabOutStore_8;
  wire[31:0] fabOutSeqClass_io_fabOutStore_7;
  wire[31:0] fabOutSeqClass_io_fabOutStore_6;
  wire[31:0] fabOutSeqClass_io_fabOutStore_5;
  wire[31:0] fabOutSeqClass_io_fabOutStore_4;
  wire[31:0] fabOutSeqClass_io_fabOutStore_3;
  wire[31:0] fabOutSeqClass_io_fabOutStore_2;
  wire[31:0] fabOutSeqClass_io_fabOutStore_1;
  wire[31:0] fabOutSeqClass_io_fabOutStore_0;
  wire fabOutSeqClass_io_fabOutStoreValid_19;
  wire fabOutSeqClass_io_fabOutStoreValid_18;
  wire fabOutSeqClass_io_fabOutStoreValid_17;
  wire fabOutSeqClass_io_fabOutStoreValid_16;
  wire fabOutSeqClass_io_fabOutStoreValid_15;
  wire fabOutSeqClass_io_fabOutStoreValid_14;
  wire fabOutSeqClass_io_fabOutStoreValid_13;
  wire fabOutSeqClass_io_fabOutStoreValid_12;
  wire fabOutSeqClass_io_fabOutStoreValid_11;
  wire fabOutSeqClass_io_fabOutStoreValid_10;
  wire fabOutSeqClass_io_fabOutStoreValid_9;
  wire fabOutSeqClass_io_fabOutStoreValid_8;
  wire fabOutSeqClass_io_fabOutStoreValid_7;
  wire fabOutSeqClass_io_fabOutStoreValid_6;
  wire fabOutSeqClass_io_fabOutStoreValid_5;
  wire fabOutSeqClass_io_fabOutStoreValid_4;
  wire fabOutSeqClass_io_fabOutStoreValid_3;
  wire fabOutSeqClass_io_fabOutStoreValid_2;
  wire fabOutSeqClass_io_fabOutStoreValid_1;
  wire fabOutSeqClass_io_fabOutStoreValid_0;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_7;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_6;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_5;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_4;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_3;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_2;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_1;
  wire[87:0] fabOutSeqClass_io_fabOutLoc_0;
  wire fabOutSeqClass_io_fabOutLocValid_7;
  wire fabOutSeqClass_io_fabOutLocValid_6;
  wire fabOutSeqClass_io_fabOutLocValid_5;
  wire fabOutSeqClass_io_fabOutLocValid_4;
  wire fabOutSeqClass_io_fabOutLocValid_3;
  wire fabOutSeqClass_io_fabOutLocValid_2;
  wire fabOutSeqClass_io_fabOutLocValid_1;
  wire fabOutSeqClass_io_fabOutLocValid_0;
  wire[31:0] fabInSeqClass_io_fabInData_19;
  wire[31:0] fabInSeqClass_io_fabInData_18;
  wire[31:0] fabInSeqClass_io_fabInData_17;
  wire[31:0] fabInSeqClass_io_fabInData_16;
  wire[31:0] fabInSeqClass_io_fabInData_15;
  wire[31:0] fabInSeqClass_io_fabInData_14;
  wire[31:0] fabInSeqClass_io_fabInData_13;
  wire[31:0] fabInSeqClass_io_fabInData_12;
  wire[31:0] fabInSeqClass_io_fabInData_11;
  wire[31:0] fabInSeqClass_io_fabInData_10;
  wire[31:0] fabInSeqClass_io_fabInData_9;
  wire[31:0] fabInSeqClass_io_fabInData_8;
  wire[31:0] fabInSeqClass_io_fabInData_7;
  wire[31:0] fabInSeqClass_io_fabInData_6;
  wire[31:0] fabInSeqClass_io_fabInData_5;
  wire[31:0] fabInSeqClass_io_fabInData_4;
  wire[31:0] fabInSeqClass_io_fabInData_3;
  wire[31:0] fabInSeqClass_io_fabInData_2;
  wire[31:0] fabInSeqClass_io_fabInData_1;
  wire[31:0] fabInSeqClass_io_fabInData_0;
  wire fabInSeqClass_io_fabInValid_19;
  wire fabInSeqClass_io_fabInValid_18;
  wire fabInSeqClass_io_fabInValid_17;
  wire fabInSeqClass_io_fabInValid_16;
  wire fabInSeqClass_io_fabInValid_15;
  wire fabInSeqClass_io_fabInValid_14;
  wire fabInSeqClass_io_fabInValid_13;
  wire fabInSeqClass_io_fabInValid_12;
  wire fabInSeqClass_io_fabInValid_11;
  wire fabInSeqClass_io_fabInValid_10;
  wire fabInSeqClass_io_fabInValid_9;
  wire fabInSeqClass_io_fabInValid_8;
  wire fabInSeqClass_io_fabInValid_7;
  wire fabInSeqClass_io_fabInValid_6;
  wire fabInSeqClass_io_fabInValid_5;
  wire fabInSeqClass_io_fabInValid_4;
  wire fabInSeqClass_io_fabInValid_3;
  wire fabInSeqClass_io_fabInValid_2;
  wire fabInSeqClass_io_fabInValid_1;
  wire fabInSeqClass_io_fabInValid_0;
  wire fabInSeqClass_io_loadStoreRdy_7;
  wire fabInSeqClass_io_loadStoreRdy_6;
  wire fabInSeqClass_io_loadStoreRdy_5;
  wire fabInSeqClass_io_loadStoreRdy_4;
  wire fabInSeqClass_io_loadStoreRdy_3;
  wire fabInSeqClass_io_loadStoreRdy_2;
  wire fabInSeqClass_io_loadStoreRdy_1;
  wire fabInSeqClass_io_loadStoreRdy_0;
  wire fabInSeqClass_io_fabStoreRdy_7;
  wire fabInSeqClass_io_fabStoreRdy_6;
  wire fabInSeqClass_io_fabStoreRdy_5;
  wire fabInSeqClass_io_fabStoreRdy_4;
  wire fabInSeqClass_io_fabStoreRdy_3;
  wire fabInSeqClass_io_fabStoreRdy_2;
  wire fabInSeqClass_io_fabStoreRdy_1;
  wire fabInSeqClass_io_fabStoreRdy_0;


  assign T0 = fabOutSeqClass_io_fabOutLoc_0[6'h25:1'h0];
  assign T1 = fabOutSeqClass_io_fabOutLoc_1[6'h25:1'h0];
  assign T2 = fabOutSeqClass_io_fabOutLoc_2[6'h25:1'h0];
  assign T3 = fabOutSeqClass_io_fabOutLoc_3[6'h25:1'h0];
  assign T4 = fabOutSeqClass_io_fabOutLoc_4[6'h25:1'h0];
  assign T5 = fabOutSeqClass_io_fabOutLoc_5[6'h25:1'h0];
  assign T6 = fabOutSeqClass_io_fabOutLoc_6[6'h25:1'h0];
  assign T7 = fabOutSeqClass_io_fabOutLoc_7[6'h25:1'h0];
  assign io_fabOutRdy_0 = fabOutSeqClass_io_fabOutRdy_0;
  assign io_fabOutRdy_1 = fabOutSeqClass_io_fabOutRdy_1;
  assign io_fabOutRdy_2 = fabOutSeqClass_io_fabOutRdy_2;
  assign io_fabOutRdy_3 = fabOutSeqClass_io_fabOutRdy_3;
  assign io_fabOutRdy_4 = fabOutSeqClass_io_fabOutRdy_4;
  assign io_fabOutRdy_5 = fabOutSeqClass_io_fabOutRdy_5;
  assign io_fabOutRdy_6 = fabOutSeqClass_io_fabOutRdy_6;
  assign io_fabOutRdy_7 = fabOutSeqClass_io_fabOutRdy_7;
  assign io_fabOutRdy_8 = fabOutSeqClass_io_fabOutRdy_8;
  assign io_fabOutRdy_9 = fabOutSeqClass_io_fabOutRdy_9;
  assign io_fabOutRdy_10 = fabOutSeqClass_io_fabOutRdy_10;
  assign io_fabOutRdy_11 = fabOutSeqClass_io_fabOutRdy_11;
  assign io_fabOutRdy_12 = fabOutSeqClass_io_fabOutRdy_12;
  assign io_fabOutRdy_13 = fabOutSeqClass_io_fabOutRdy_13;
  assign io_fabOutRdy_14 = fabOutSeqClass_io_fabOutRdy_14;
  assign io_fabOutRdy_15 = fabOutSeqClass_io_fabOutRdy_15;
  assign io_fabOutRdy_16 = fabOutSeqClass_io_fabOutRdy_16;
  assign io_fabOutRdy_17 = fabOutSeqClass_io_fabOutRdy_17;
  assign io_fabOutRdy_18 = fabOutSeqClass_io_fabOutRdy_18;
  assign io_fabOutRdy_19 = fabOutSeqClass_io_fabOutRdy_19;
  assign io_fabInValid_0 = fabInSeqClass_io_fabInValid_0;
  assign io_fabInValid_1 = fabInSeqClass_io_fabInValid_1;
  assign io_fabInValid_2 = fabInSeqClass_io_fabInValid_2;
  assign io_fabInValid_3 = fabInSeqClass_io_fabInValid_3;
  assign io_fabInValid_4 = fabInSeqClass_io_fabInValid_4;
  assign io_fabInValid_5 = fabInSeqClass_io_fabInValid_5;
  assign io_fabInValid_6 = fabInSeqClass_io_fabInValid_6;
  assign io_fabInValid_7 = fabInSeqClass_io_fabInValid_7;
  assign io_fabInValid_8 = fabInSeqClass_io_fabInValid_8;
  assign io_fabInValid_9 = fabInSeqClass_io_fabInValid_9;
  assign io_fabInValid_10 = fabInSeqClass_io_fabInValid_10;
  assign io_fabInValid_11 = fabInSeqClass_io_fabInValid_11;
  assign io_fabInValid_12 = fabInSeqClass_io_fabInValid_12;
  assign io_fabInValid_13 = fabInSeqClass_io_fabInValid_13;
  assign io_fabInValid_14 = fabInSeqClass_io_fabInValid_14;
  assign io_fabInValid_15 = fabInSeqClass_io_fabInValid_15;
  assign io_fabInValid_16 = fabInSeqClass_io_fabInValid_16;
  assign io_fabInValid_17 = fabInSeqClass_io_fabInValid_17;
  assign io_fabInValid_18 = fabInSeqClass_io_fabInValid_18;
  assign io_fabInValid_19 = fabInSeqClass_io_fabInValid_19;
  assign io_fabInData_0 = fabInSeqClass_io_fabInData_0;
  assign io_fabInData_1 = fabInSeqClass_io_fabInData_1;
  assign io_fabInData_2 = fabInSeqClass_io_fabInData_2;
  assign io_fabInData_3 = fabInSeqClass_io_fabInData_3;
  assign io_fabInData_4 = fabInSeqClass_io_fabInData_4;
  assign io_fabInData_5 = fabInSeqClass_io_fabInData_5;
  assign io_fabInData_6 = fabInSeqClass_io_fabInData_6;
  assign io_fabInData_7 = fabInSeqClass_io_fabInData_7;
  assign io_fabInData_8 = fabInSeqClass_io_fabInData_8;
  assign io_fabInData_9 = fabInSeqClass_io_fabInData_9;
  assign io_fabInData_10 = fabInSeqClass_io_fabInData_10;
  assign io_fabInData_11 = fabInSeqClass_io_fabInData_11;
  assign io_fabInData_12 = fabInSeqClass_io_fabInData_12;
  assign io_fabInData_13 = fabInSeqClass_io_fabInData_13;
  assign io_fabInData_14 = fabInSeqClass_io_fabInData_14;
  assign io_fabInData_15 = fabInSeqClass_io_fabInData_15;
  assign io_fabInData_16 = fabInSeqClass_io_fabInData_16;
  assign io_fabInData_17 = fabInSeqClass_io_fabInData_17;
  assign io_fabInData_18 = fabInSeqClass_io_fabInData_18;
  assign io_fabInData_19 = fabInSeqClass_io_fabInData_19;
  assign io_storeMemValid = storeSeqClass_io_storeMemValid;
  assign io_storeMemData = storeSeqClass_io_storeMemData;
  assign io_loadRespRdy = loadSeqClass_io_loadRespRdy;
  assign io_loadRqstValid = loadSeqClass_io_loadRqstValid;
  assign io_loadRqst = loadSeqClass_io_loadRqst;
  fabInSeq fabInSeqClass(.clk(clk), .reset(reset),
       .io_inConfig( mainConfigClass_io_fabInConfig ),
       .io_inValid( mainConfigClass_io_fabInConfigValid ),
       .io_fabInData_19( fabInSeqClass_io_fabInData_19 ),
       .io_fabInData_18( fabInSeqClass_io_fabInData_18 ),
       .io_fabInData_17( fabInSeqClass_io_fabInData_17 ),
       .io_fabInData_16( fabInSeqClass_io_fabInData_16 ),
       .io_fabInData_15( fabInSeqClass_io_fabInData_15 ),
       .io_fabInData_14( fabInSeqClass_io_fabInData_14 ),
       .io_fabInData_13( fabInSeqClass_io_fabInData_13 ),
       .io_fabInData_12( fabInSeqClass_io_fabInData_12 ),
       .io_fabInData_11( fabInSeqClass_io_fabInData_11 ),
       .io_fabInData_10( fabInSeqClass_io_fabInData_10 ),
       .io_fabInData_9( fabInSeqClass_io_fabInData_9 ),
       .io_fabInData_8( fabInSeqClass_io_fabInData_8 ),
       .io_fabInData_7( fabInSeqClass_io_fabInData_7 ),
       .io_fabInData_6( fabInSeqClass_io_fabInData_6 ),
       .io_fabInData_5( fabInSeqClass_io_fabInData_5 ),
       .io_fabInData_4( fabInSeqClass_io_fabInData_4 ),
       .io_fabInData_3( fabInSeqClass_io_fabInData_3 ),
       .io_fabInData_2( fabInSeqClass_io_fabInData_2 ),
       .io_fabInData_1( fabInSeqClass_io_fabInData_1 ),
       .io_fabInData_0( fabInSeqClass_io_fabInData_0 ),
       .io_fabInValid_19( fabInSeqClass_io_fabInValid_19 ),
       .io_fabInValid_18( fabInSeqClass_io_fabInValid_18 ),
       .io_fabInValid_17( fabInSeqClass_io_fabInValid_17 ),
       .io_fabInValid_16( fabInSeqClass_io_fabInValid_16 ),
       .io_fabInValid_15( fabInSeqClass_io_fabInValid_15 ),
       .io_fabInValid_14( fabInSeqClass_io_fabInValid_14 ),
       .io_fabInValid_13( fabInSeqClass_io_fabInValid_13 ),
       .io_fabInValid_12( fabInSeqClass_io_fabInValid_12 ),
       .io_fabInValid_11( fabInSeqClass_io_fabInValid_11 ),
       .io_fabInValid_10( fabInSeqClass_io_fabInValid_10 ),
       .io_fabInValid_9( fabInSeqClass_io_fabInValid_9 ),
       .io_fabInValid_8( fabInSeqClass_io_fabInValid_8 ),
       .io_fabInValid_7( fabInSeqClass_io_fabInValid_7 ),
       .io_fabInValid_6( fabInSeqClass_io_fabInValid_6 ),
       .io_fabInValid_5( fabInSeqClass_io_fabInValid_5 ),
       .io_fabInValid_4( fabInSeqClass_io_fabInValid_4 ),
       .io_fabInValid_3( fabInSeqClass_io_fabInValid_3 ),
       .io_fabInValid_2( fabInSeqClass_io_fabInValid_2 ),
       .io_fabInValid_1( fabInSeqClass_io_fabInValid_1 ),
       .io_fabInValid_0( fabInSeqClass_io_fabInValid_0 ),
       .io_fabInRdy_19( io_fabInRdy_19 ),
       .io_fabInRdy_18( io_fabInRdy_18 ),
       .io_fabInRdy_17( io_fabInRdy_17 ),
       .io_fabInRdy_16( io_fabInRdy_16 ),
       .io_fabInRdy_15( io_fabInRdy_15 ),
       .io_fabInRdy_14( io_fabInRdy_14 ),
       .io_fabInRdy_13( io_fabInRdy_13 ),
       .io_fabInRdy_12( io_fabInRdy_12 ),
       .io_fabInRdy_11( io_fabInRdy_11 ),
       .io_fabInRdy_10( io_fabInRdy_10 ),
       .io_fabInRdy_9( io_fabInRdy_9 ),
       .io_fabInRdy_8( io_fabInRdy_8 ),
       .io_fabInRdy_7( io_fabInRdy_7 ),
       .io_fabInRdy_6( io_fabInRdy_6 ),
       .io_fabInRdy_5( io_fabInRdy_5 ),
       .io_fabInRdy_4( io_fabInRdy_4 ),
       .io_fabInRdy_3( io_fabInRdy_3 ),
       .io_fabInRdy_2( io_fabInRdy_2 ),
       .io_fabInRdy_1( io_fabInRdy_1 ),
       .io_fabInRdy_0( io_fabInRdy_0 ),
       .io_loadStore_7( loadSeqClass_io_memBankEnq_7 ),
       .io_loadStore_6( loadSeqClass_io_memBankEnq_6 ),
       .io_loadStore_5( loadSeqClass_io_memBankEnq_5 ),
       .io_loadStore_4( loadSeqClass_io_memBankEnq_4 ),
       .io_loadStore_3( loadSeqClass_io_memBankEnq_3 ),
       .io_loadStore_2( loadSeqClass_io_memBankEnq_2 ),
       .io_loadStore_1( loadSeqClass_io_memBankEnq_1 ),
       .io_loadStore_0( loadSeqClass_io_memBankEnq_0 ),
       .io_loadStoreValid_7( loadSeqClass_io_memBankValid_7 ),
       .io_loadStoreValid_6( loadSeqClass_io_memBankValid_6 ),
       .io_loadStoreValid_5( loadSeqClass_io_memBankValid_5 ),
       .io_loadStoreValid_4( loadSeqClass_io_memBankValid_4 ),
       .io_loadStoreValid_3( loadSeqClass_io_memBankValid_3 ),
       .io_loadStoreValid_2( loadSeqClass_io_memBankValid_2 ),
       .io_loadStoreValid_1( loadSeqClass_io_memBankValid_1 ),
       .io_loadStoreValid_0( loadSeqClass_io_memBankValid_0 ),
       .io_loadStoreRdy_7( fabInSeqClass_io_loadStoreRdy_7 ),
       .io_loadStoreRdy_6( fabInSeqClass_io_loadStoreRdy_6 ),
       .io_loadStoreRdy_5( fabInSeqClass_io_loadStoreRdy_5 ),
       .io_loadStoreRdy_4( fabInSeqClass_io_loadStoreRdy_4 ),
       .io_loadStoreRdy_3( fabInSeqClass_io_loadStoreRdy_3 ),
       .io_loadStoreRdy_2( fabInSeqClass_io_loadStoreRdy_2 ),
       .io_loadStoreRdy_1( fabInSeqClass_io_loadStoreRdy_1 ),
       .io_loadStoreRdy_0( fabInSeqClass_io_loadStoreRdy_0 ),
       .io_fabStore_7( T7 ),
       .io_fabStore_6( T6 ),
       .io_fabStore_5( T5 ),
       .io_fabStore_4( T4 ),
       .io_fabStore_3( T3 ),
       .io_fabStore_2( T2 ),
       .io_fabStore_1( T1 ),
       .io_fabStore_0( T0 ),
       .io_fabStoreValid_7( fabOutSeqClass_io_fabOutLocValid_7 ),
       .io_fabStoreValid_6( fabOutSeqClass_io_fabOutLocValid_6 ),
       .io_fabStoreValid_5( fabOutSeqClass_io_fabOutLocValid_5 ),
       .io_fabStoreValid_4( fabOutSeqClass_io_fabOutLocValid_4 ),
       .io_fabStoreValid_3( fabOutSeqClass_io_fabOutLocValid_3 ),
       .io_fabStoreValid_2( fabOutSeqClass_io_fabOutLocValid_2 ),
       .io_fabStoreValid_1( fabOutSeqClass_io_fabOutLocValid_1 ),
       .io_fabStoreValid_0( fabOutSeqClass_io_fabOutLocValid_0 ),
       .io_fabStoreRdy_7( fabInSeqClass_io_fabStoreRdy_7 ),
       .io_fabStoreRdy_6( fabInSeqClass_io_fabStoreRdy_6 ),
       .io_fabStoreRdy_5( fabInSeqClass_io_fabStoreRdy_5 ),
       .io_fabStoreRdy_4( fabInSeqClass_io_fabStoreRdy_4 ),
       .io_fabStoreRdy_3( fabInSeqClass_io_fabStoreRdy_3 ),
       .io_fabStoreRdy_2( fabInSeqClass_io_fabStoreRdy_2 ),
       .io_fabStoreRdy_1( fabInSeqClass_io_fabStoreRdy_1 ),
       .io_fabStoreRdy_0( fabInSeqClass_io_fabStoreRdy_0 )
       //.io_computeDone(  )
  );
  fabOutSeqTop fabOutSeqClass(.clk(clk), .reset(reset),
       .io_inConfig( mainConfigClass_io_fabOutConfig ),
       .io_inValid( mainConfigClass_io_fabOutConfigValid ),
       .io_fabOut_19( io_fabOut_19 ),
       .io_fabOut_18( io_fabOut_18 ),
       .io_fabOut_17( io_fabOut_17 ),
       .io_fabOut_16( io_fabOut_16 ),
       .io_fabOut_15( io_fabOut_15 ),
       .io_fabOut_14( io_fabOut_14 ),
       .io_fabOut_13( io_fabOut_13 ),
       .io_fabOut_12( io_fabOut_12 ),
       .io_fabOut_11( io_fabOut_11 ),
       .io_fabOut_10( io_fabOut_10 ),
       .io_fabOut_9( io_fabOut_9 ),
       .io_fabOut_8( io_fabOut_8 ),
       .io_fabOut_7( io_fabOut_7 ),
       .io_fabOut_6( io_fabOut_6 ),
       .io_fabOut_5( io_fabOut_5 ),
       .io_fabOut_4( io_fabOut_4 ),
       .io_fabOut_3( io_fabOut_3 ),
       .io_fabOut_2( io_fabOut_2 ),
       .io_fabOut_1( io_fabOut_1 ),
       .io_fabOut_0( io_fabOut_0 ),
       .io_fabOutValid_19( io_fabOutValid_19 ),
       .io_fabOutValid_18( io_fabOutValid_18 ),
       .io_fabOutValid_17( io_fabOutValid_17 ),
       .io_fabOutValid_16( io_fabOutValid_16 ),
       .io_fabOutValid_15( io_fabOutValid_15 ),
       .io_fabOutValid_14( io_fabOutValid_14 ),
       .io_fabOutValid_13( io_fabOutValid_13 ),
       .io_fabOutValid_12( io_fabOutValid_12 ),
       .io_fabOutValid_11( io_fabOutValid_11 ),
       .io_fabOutValid_10( io_fabOutValid_10 ),
       .io_fabOutValid_9( io_fabOutValid_9 ),
       .io_fabOutValid_8( io_fabOutValid_8 ),
       .io_fabOutValid_7( io_fabOutValid_7 ),
       .io_fabOutValid_6( io_fabOutValid_6 ),
       .io_fabOutValid_5( io_fabOutValid_5 ),
       .io_fabOutValid_4( io_fabOutValid_4 ),
       .io_fabOutValid_3( io_fabOutValid_3 ),
       .io_fabOutValid_2( io_fabOutValid_2 ),
       .io_fabOutValid_1( io_fabOutValid_1 ),
       .io_fabOutValid_0( io_fabOutValid_0 ),
       .io_fabOutRdy_19( fabOutSeqClass_io_fabOutRdy_19 ),
       .io_fabOutRdy_18( fabOutSeqClass_io_fabOutRdy_18 ),
       .io_fabOutRdy_17( fabOutSeqClass_io_fabOutRdy_17 ),
       .io_fabOutRdy_16( fabOutSeqClass_io_fabOutRdy_16 ),
       .io_fabOutRdy_15( fabOutSeqClass_io_fabOutRdy_15 ),
       .io_fabOutRdy_14( fabOutSeqClass_io_fabOutRdy_14 ),
       .io_fabOutRdy_13( fabOutSeqClass_io_fabOutRdy_13 ),
       .io_fabOutRdy_12( fabOutSeqClass_io_fabOutRdy_12 ),
       .io_fabOutRdy_11( fabOutSeqClass_io_fabOutRdy_11 ),
       .io_fabOutRdy_10( fabOutSeqClass_io_fabOutRdy_10 ),
       .io_fabOutRdy_9( fabOutSeqClass_io_fabOutRdy_9 ),
       .io_fabOutRdy_8( fabOutSeqClass_io_fabOutRdy_8 ),
       .io_fabOutRdy_7( fabOutSeqClass_io_fabOutRdy_7 ),
       .io_fabOutRdy_6( fabOutSeqClass_io_fabOutRdy_6 ),
       .io_fabOutRdy_5( fabOutSeqClass_io_fabOutRdy_5 ),
       .io_fabOutRdy_4( fabOutSeqClass_io_fabOutRdy_4 ),
       .io_fabOutRdy_3( fabOutSeqClass_io_fabOutRdy_3 ),
       .io_fabOutRdy_2( fabOutSeqClass_io_fabOutRdy_2 ),
       .io_fabOutRdy_1( fabOutSeqClass_io_fabOutRdy_1 ),
       .io_fabOutRdy_0( fabOutSeqClass_io_fabOutRdy_0 ),
       .io_fabOutStore_19( fabOutSeqClass_io_fabOutStore_19 ),
       .io_fabOutStore_18( fabOutSeqClass_io_fabOutStore_18 ),
       .io_fabOutStore_17( fabOutSeqClass_io_fabOutStore_17 ),
       .io_fabOutStore_16( fabOutSeqClass_io_fabOutStore_16 ),
       .io_fabOutStore_15( fabOutSeqClass_io_fabOutStore_15 ),
       .io_fabOutStore_14( fabOutSeqClass_io_fabOutStore_14 ),
       .io_fabOutStore_13( fabOutSeqClass_io_fabOutStore_13 ),
       .io_fabOutStore_12( fabOutSeqClass_io_fabOutStore_12 ),
       .io_fabOutStore_11( fabOutSeqClass_io_fabOutStore_11 ),
       .io_fabOutStore_10( fabOutSeqClass_io_fabOutStore_10 ),
       .io_fabOutStore_9( fabOutSeqClass_io_fabOutStore_9 ),
       .io_fabOutStore_8( fabOutSeqClass_io_fabOutStore_8 ),
       .io_fabOutStore_7( fabOutSeqClass_io_fabOutStore_7 ),
       .io_fabOutStore_6( fabOutSeqClass_io_fabOutStore_6 ),
       .io_fabOutStore_5( fabOutSeqClass_io_fabOutStore_5 ),
       .io_fabOutStore_4( fabOutSeqClass_io_fabOutStore_4 ),
       .io_fabOutStore_3( fabOutSeqClass_io_fabOutStore_3 ),
       .io_fabOutStore_2( fabOutSeqClass_io_fabOutStore_2 ),
       .io_fabOutStore_1( fabOutSeqClass_io_fabOutStore_1 ),
       .io_fabOutStore_0( fabOutSeqClass_io_fabOutStore_0 ),
       .io_fabOutStoreValid_19( fabOutSeqClass_io_fabOutStoreValid_19 ),
       .io_fabOutStoreValid_18( fabOutSeqClass_io_fabOutStoreValid_18 ),
       .io_fabOutStoreValid_17( fabOutSeqClass_io_fabOutStoreValid_17 ),
       .io_fabOutStoreValid_16( fabOutSeqClass_io_fabOutStoreValid_16 ),
       .io_fabOutStoreValid_15( fabOutSeqClass_io_fabOutStoreValid_15 ),
       .io_fabOutStoreValid_14( fabOutSeqClass_io_fabOutStoreValid_14 ),
       .io_fabOutStoreValid_13( fabOutSeqClass_io_fabOutStoreValid_13 ),
       .io_fabOutStoreValid_12( fabOutSeqClass_io_fabOutStoreValid_12 ),
       .io_fabOutStoreValid_11( fabOutSeqClass_io_fabOutStoreValid_11 ),
       .io_fabOutStoreValid_10( fabOutSeqClass_io_fabOutStoreValid_10 ),
       .io_fabOutStoreValid_9( fabOutSeqClass_io_fabOutStoreValid_9 ),
       .io_fabOutStoreValid_8( fabOutSeqClass_io_fabOutStoreValid_8 ),
       .io_fabOutStoreValid_7( fabOutSeqClass_io_fabOutStoreValid_7 ),
       .io_fabOutStoreValid_6( fabOutSeqClass_io_fabOutStoreValid_6 ),
       .io_fabOutStoreValid_5( fabOutSeqClass_io_fabOutStoreValid_5 ),
       .io_fabOutStoreValid_4( fabOutSeqClass_io_fabOutStoreValid_4 ),
       .io_fabOutStoreValid_3( fabOutSeqClass_io_fabOutStoreValid_3 ),
       .io_fabOutStoreValid_2( fabOutSeqClass_io_fabOutStoreValid_2 ),
       .io_fabOutStoreValid_1( fabOutSeqClass_io_fabOutStoreValid_1 ),
       .io_fabOutStoreValid_0( fabOutSeqClass_io_fabOutStoreValid_0 ),
       //.io_fabOutStoreRdy_19(  )
       //.io_fabOutStoreRdy_18(  )
       //.io_fabOutStoreRdy_17(  )
       //.io_fabOutStoreRdy_16(  )
       //.io_fabOutStoreRdy_15(  )
       //.io_fabOutStoreRdy_14(  )
       //.io_fabOutStoreRdy_13(  )
       //.io_fabOutStoreRdy_12(  )
       //.io_fabOutStoreRdy_11(  )
       //.io_fabOutStoreRdy_10(  )
       //.io_fabOutStoreRdy_9(  )
       //.io_fabOutStoreRdy_8(  )
       //.io_fabOutStoreRdy_7(  )
       //.io_fabOutStoreRdy_6(  )
       //.io_fabOutStoreRdy_5(  )
       //.io_fabOutStoreRdy_4(  )
       //.io_fabOutStoreRdy_3(  )
       //.io_fabOutStoreRdy_2(  )
       //.io_fabOutStoreRdy_1(  )
       //.io_fabOutStoreRdy_0(  )
       .io_fabOutLoc_7( fabOutSeqClass_io_fabOutLoc_7 ),
       .io_fabOutLoc_6( fabOutSeqClass_io_fabOutLoc_6 ),
       .io_fabOutLoc_5( fabOutSeqClass_io_fabOutLoc_5 ),
       .io_fabOutLoc_4( fabOutSeqClass_io_fabOutLoc_4 ),
       .io_fabOutLoc_3( fabOutSeqClass_io_fabOutLoc_3 ),
       .io_fabOutLoc_2( fabOutSeqClass_io_fabOutLoc_2 ),
       .io_fabOutLoc_1( fabOutSeqClass_io_fabOutLoc_1 ),
       .io_fabOutLoc_0( fabOutSeqClass_io_fabOutLoc_0 ),
       .io_fabOutLocValid_7( fabOutSeqClass_io_fabOutLocValid_7 ),
       .io_fabOutLocValid_6( fabOutSeqClass_io_fabOutLocValid_6 ),
       .io_fabOutLocValid_5( fabOutSeqClass_io_fabOutLocValid_5 ),
       .io_fabOutLocValid_4( fabOutSeqClass_io_fabOutLocValid_4 ),
       .io_fabOutLocValid_3( fabOutSeqClass_io_fabOutLocValid_3 ),
       .io_fabOutLocValid_2( fabOutSeqClass_io_fabOutLocValid_2 ),
       .io_fabOutLocValid_1( fabOutSeqClass_io_fabOutLocValid_1 ),
       .io_fabOutLocValid_0( fabOutSeqClass_io_fabOutLocValid_0 ),
       .io_fabOutLocRdy_7( fabInSeqClass_io_fabStoreRdy_7 ),
       .io_fabOutLocRdy_6( fabInSeqClass_io_fabStoreRdy_6 ),
       .io_fabOutLocRdy_5( fabInSeqClass_io_fabStoreRdy_5 ),
       .io_fabOutLocRdy_4( fabInSeqClass_io_fabStoreRdy_4 ),
       .io_fabOutLocRdy_3( fabInSeqClass_io_fabStoreRdy_3 ),
       .io_fabOutLocRdy_2( fabInSeqClass_io_fabStoreRdy_2 ),
       .io_fabOutLocRdy_1( fabInSeqClass_io_fabStoreRdy_1 ),
       .io_fabOutLocRdy_0( fabInSeqClass_io_fabStoreRdy_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabOutSeqClass.io_fabOutStoreRdy_19 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_18 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_17 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_16 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_15 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_14 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_13 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_12 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_11 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_10 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_9 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_8 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_7 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_6 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_5 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_4 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_3 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_2 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_1 = {1{$random}};
    assign fabOutSeqClass.io_fabOutStoreRdy_0 = {1{$random}};
// synthesis translate_on
`endif
  loadSeq loadSeqClass(.clk(clk), .reset(reset),
       .io_inConfig( mainConfigClass_io_loadConfig ),
       .io_inValid( mainConfigClass_io_loadConfigValid ),
       .io_loadRqst( loadSeqClass_io_loadRqst ),
       .io_loadRqstValid( loadSeqClass_io_loadRqstValid ),
       .io_loadRqstRdy( io_loadRqstRdy ),
       .io_loadResp( io_loadResp ),
       .io_loadRespValid( io_loadRespValid ),
       .io_loadRespRdy( loadSeqClass_io_loadRespRdy ),
       .io_memBankEnq_7( loadSeqClass_io_memBankEnq_7 ),
       .io_memBankEnq_6( loadSeqClass_io_memBankEnq_6 ),
       .io_memBankEnq_5( loadSeqClass_io_memBankEnq_5 ),
       .io_memBankEnq_4( loadSeqClass_io_memBankEnq_4 ),
       .io_memBankEnq_3( loadSeqClass_io_memBankEnq_3 ),
       .io_memBankEnq_2( loadSeqClass_io_memBankEnq_2 ),
       .io_memBankEnq_1( loadSeqClass_io_memBankEnq_1 ),
       .io_memBankEnq_0( loadSeqClass_io_memBankEnq_0 ),
       .io_memBankValid_7( loadSeqClass_io_memBankValid_7 ),
       .io_memBankValid_6( loadSeqClass_io_memBankValid_6 ),
       .io_memBankValid_5( loadSeqClass_io_memBankValid_5 ),
       .io_memBankValid_4( loadSeqClass_io_memBankValid_4 ),
       .io_memBankValid_3( loadSeqClass_io_memBankValid_3 ),
       .io_memBankValid_2( loadSeqClass_io_memBankValid_2 ),
       .io_memBankValid_1( loadSeqClass_io_memBankValid_1 ),
       .io_memBankValid_0( loadSeqClass_io_memBankValid_0 ),
       .io_memBankRdy_7( fabInSeqClass_io_loadStoreRdy_7 ),
       .io_memBankRdy_6( fabInSeqClass_io_loadStoreRdy_6 ),
       .io_memBankRdy_5( fabInSeqClass_io_loadStoreRdy_5 ),
       .io_memBankRdy_4( fabInSeqClass_io_loadStoreRdy_4 ),
       .io_memBankRdy_3( fabInSeqClass_io_loadStoreRdy_3 ),
       .io_memBankRdy_2( fabInSeqClass_io_loadStoreRdy_2 ),
       .io_memBankRdy_1( fabInSeqClass_io_loadStoreRdy_1 ),
       .io_memBankRdy_0( fabInSeqClass_io_loadStoreRdy_0 )
  );
  storeSeq storeSeqClass(.clk(clk), .reset(reset),
       .io_inConfig( mainConfigClass_io_storeConfig ),
       .io_inValid( mainConfigClass_io_storeConfigValid ),
       .io_fabOutToStore_19( fabOutSeqClass_io_fabOutStore_19 ),
       .io_fabOutToStore_18( fabOutSeqClass_io_fabOutStore_18 ),
       .io_fabOutToStore_17( fabOutSeqClass_io_fabOutStore_17 ),
       .io_fabOutToStore_16( fabOutSeqClass_io_fabOutStore_16 ),
       .io_fabOutToStore_15( fabOutSeqClass_io_fabOutStore_15 ),
       .io_fabOutToStore_14( fabOutSeqClass_io_fabOutStore_14 ),
       .io_fabOutToStore_13( fabOutSeqClass_io_fabOutStore_13 ),
       .io_fabOutToStore_12( fabOutSeqClass_io_fabOutStore_12 ),
       .io_fabOutToStore_11( fabOutSeqClass_io_fabOutStore_11 ),
       .io_fabOutToStore_10( fabOutSeqClass_io_fabOutStore_10 ),
       .io_fabOutToStore_9( fabOutSeqClass_io_fabOutStore_9 ),
       .io_fabOutToStore_8( fabOutSeqClass_io_fabOutStore_8 ),
       .io_fabOutToStore_7( fabOutSeqClass_io_fabOutStore_7 ),
       .io_fabOutToStore_6( fabOutSeqClass_io_fabOutStore_6 ),
       .io_fabOutToStore_5( fabOutSeqClass_io_fabOutStore_5 ),
       .io_fabOutToStore_4( fabOutSeqClass_io_fabOutStore_4 ),
       .io_fabOutToStore_3( fabOutSeqClass_io_fabOutStore_3 ),
       .io_fabOutToStore_2( fabOutSeqClass_io_fabOutStore_2 ),
       .io_fabOutToStore_1( fabOutSeqClass_io_fabOutStore_1 ),
       .io_fabOutToStore_0( fabOutSeqClass_io_fabOutStore_0 ),
       .io_fabOutToStoreValid_19( fabOutSeqClass_io_fabOutStoreValid_19 ),
       .io_fabOutToStoreValid_18( fabOutSeqClass_io_fabOutStoreValid_18 ),
       .io_fabOutToStoreValid_17( fabOutSeqClass_io_fabOutStoreValid_17 ),
       .io_fabOutToStoreValid_16( fabOutSeqClass_io_fabOutStoreValid_16 ),
       .io_fabOutToStoreValid_15( fabOutSeqClass_io_fabOutStoreValid_15 ),
       .io_fabOutToStoreValid_14( fabOutSeqClass_io_fabOutStoreValid_14 ),
       .io_fabOutToStoreValid_13( fabOutSeqClass_io_fabOutStoreValid_13 ),
       .io_fabOutToStoreValid_12( fabOutSeqClass_io_fabOutStoreValid_12 ),
       .io_fabOutToStoreValid_11( fabOutSeqClass_io_fabOutStoreValid_11 ),
       .io_fabOutToStoreValid_10( fabOutSeqClass_io_fabOutStoreValid_10 ),
       .io_fabOutToStoreValid_9( fabOutSeqClass_io_fabOutStoreValid_9 ),
       .io_fabOutToStoreValid_8( fabOutSeqClass_io_fabOutStoreValid_8 ),
       .io_fabOutToStoreValid_7( fabOutSeqClass_io_fabOutStoreValid_7 ),
       .io_fabOutToStoreValid_6( fabOutSeqClass_io_fabOutStoreValid_6 ),
       .io_fabOutToStoreValid_5( fabOutSeqClass_io_fabOutStoreValid_5 ),
       .io_fabOutToStoreValid_4( fabOutSeqClass_io_fabOutStoreValid_4 ),
       .io_fabOutToStoreValid_3( fabOutSeqClass_io_fabOutStoreValid_3 ),
       .io_fabOutToStoreValid_2( fabOutSeqClass_io_fabOutStoreValid_2 ),
       .io_fabOutToStoreValid_1( fabOutSeqClass_io_fabOutStoreValid_1 ),
       .io_fabOutToStoreValid_0( fabOutSeqClass_io_fabOutStoreValid_0 ),
       .io_storeMemData( storeSeqClass_io_storeMemData ),
       .io_storeMemValid( storeSeqClass_io_storeMemValid ),
       .io_storeMemRdy( io_storeMemRdy )
       //.io_computeDone(  )
  );
  mainConfigure mainConfigClass(.clk(clk), .reset(reset),
       .io_configData( io_inConfig ),
       .io_configDataValid( io_inValid ),
       .io_loadConfig( mainConfigClass_io_loadConfig ),
       .io_loadConfigValid( mainConfigClass_io_loadConfigValid ),
       .io_storeConfig( mainConfigClass_io_storeConfig ),
       .io_storeConfigValid( mainConfigClass_io_storeConfigValid ),
       .io_fabInConfig( mainConfigClass_io_fabInConfig ),
       .io_fabInConfigValid( mainConfigClass_io_fabInConfigValid ),
       .io_fabOutConfig( mainConfigClass_io_fabOutConfig ),
       .io_fabOutConfigValid( mainConfigClass_io_fabOutConfigValid )
       //.io_fabConfig(  )
       //.io_fabConfigValid(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign mainConfigClass.io_loadConfig = {1{$random}};
    assign mainConfigClass.io_loadConfigValid = {1{$random}};
// synthesis translate_on
`endif
  fabricConfigureTop fabConfigClass(.clk(clk), .reset(reset),
       //.io_inConfig(  )
       //.io_outConfig_5(  )
       //.io_outConfig_4(  )
       //.io_outConfig_3(  )
       //.io_outConfig_2(  )
       //.io_outConfig_1(  )
       //.io_outConfig_0(  )
       //.io_rst(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign fabConfigClass.io_inConfig = {1{$random}};
    assign fabConfigClass.io_rst = {1{$random}};
// synthesis translate_on
`endif
endmodule

